module RocketTile
   (O,
    mem_reg_replay_reg,
    ADDRARDADDR,
    ADDRBWRADDR,
    sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_opcode,
    sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_param,
    sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_size,
    sbus_auto_coupler_to_mbus_nodelay_out_c_bits_size,
    DOA,
    \remainder_reg[107] ,
    \remainder_reg[111] ,
    \remainder_reg[115] ,
    \remainder_reg[115]_0 ,
    \remainder_reg[103] ,
    \remainder_reg[107]_0 ,
    \remainder_reg[111]_0 ,
    \remainder_reg[115]_1 ,
    data_arrays_0_0_reg_i_52,
    sbus_auto_coupler_from_tile_named_tile_fixer_in_d_ready,
    tag_array_0_reg_i_13__0,
    s2_valid_reg,
    D,
    \_T_767_reg[2] ,
    \_T_5874_reg[1] ,
    sbus_auto_coupler_from_tile_named_tile_fixer_in_a_valid,
    \_T_5874_reg[0] ,
    ram_address__T_63_data,
    count_reg,
    _T_1053_reg,
    got_e_reg,
    got_e_reg_0,
    Q,
    \_T_5369_reg[5] ,
    \_T_6233_reg[5] ,
    \_T_6215_reg[3] ,
    \_T_6215_reg[2] ,
    \_T_6215_reg[1] ,
    \_T_5856_reg[0] ,
    \_T_5351_reg[0] ,
    \_T_5351_reg[3] ,
    \_T_5856_reg[3] ,
    DIB,
    \ram_opcode_reg[1] ,
    \saved_address_reg[1] ,
    \_T_6233_reg[0] ,
    \saved_address_reg[1]_0 ,
    \saved_address_reg[7] ,
    \saved_address_reg[7]_0 ,
    \saved_address_reg[7]_1 ,
    \saved_address_reg[7]_2 ,
    \saved_address_reg[7]_3 ,
    \saved_address_reg[7]_4 ,
    system_bus_xbar_auto_out_3_a_bits_param,
    DIA,
    \_T_6233_reg[1] ,
    \_T_4992_reg[2] ,
    \_T_5874_reg[2] ,
    \_T_6233_reg[0]_0 ,
    _T_5195_0_reg,
    value_1_reg,
    \_T_4992_reg[3] ,
    \_T_5856_reg[5] ,
    \_T_4992_reg[7] ,
    \_T_4992_reg[6] ,
    \_T_4992_reg[8] ,
    \_T_5856_reg[1] ,
    \_T_5856_reg[2] ,
    maybe_full_reg,
    \_T_1057_reg[1] ,
    \_T_1057_reg[0] ,
    \_T_1057_reg[1]_0 ,
    \_T_1057_reg[0]_0 ,
    \ram_strb_reg[0] ,
    _T_920_0_reg,
    \ram_strb_reg[2] ,
    \ram_strb_reg[4] ,
    \ram_strb_reg[0]_0 ,
    \ram_strb_reg[2]_0 ,
    \ram_strb_reg[4]_0 ,
    \ram_strb_reg[6] ,
    \ram_strb_reg[6]_0 ,
    \ram_strb_reg[1] ,
    \ram_strb_reg[3] ,
    \ram_strb_reg[5] ,
    \ram_strb_reg[7] ,
    \ram_id_reg[4] ,
    \ram_id_reg[0] ,
    ram_source__T_63_data,
    \ram_id_reg[3] ,
    \ram_id_reg[5] ,
    \ram_user_reg[6] ,
    _T_940_0,
    _T_920_3_reg,
    maybe_full_reg_0,
    \value_1_reg[1] ,
    \value_1_reg[0] ,
    _T_1670_reg,
    _T_642_1_reg,
    count_reg_0,
    count_reg_1,
    count_reg_2,
    count_reg_3,
    count_reg_4,
    count_reg_5,
    count_reg_6,
    \source_reg[1] ,
    ram_mask__T_63_data,
    ram_data__T_63_data,
    \ram_data_reg[63] ,
    _GEN_61,
    _GEN_55,
    host_clk,
    target_reset,
    sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_opcode,
    sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_size,
    sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_sink,
    sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_error,
    tile_auto_int_sync_xing_sinklzy_in_2_sync_0,
    S,
    \remainder_reg[64] ,
    \remainder_reg[64]_0 ,
    \remainder_reg[64]_1 ,
    DI,
    data_arrays_0_0_reg_i_44,
    data_arrays_0_0_reg_i_45,
    data_arrays_0_0_reg_i_46,
    data_arrays_0_0_reg_i_47,
    data_arrays_0_0_reg_i_48,
    data_arrays_0_0_reg_i_49,
    data_arrays_0_0_reg_i_50,
    data_arrays_0_0_reg_i_51,
    data_arrays_0_0_reg_i_52_0,
    sbus_auto_coupler_from_tile_named_tile_fixer_in_b_valid,
    sbus_auto_coupler_from_tile_named_tile_fixer_in_a_ready,
    data_arrays_1_0_reg_i_11,
    data_arrays_1_0_reg_i_12,
    data_arrays_1_0_reg_i_13,
    data_arrays_1_0_reg_i_14,
    data_arrays_1_0_reg_i_15,
    data_arrays_1_0_reg_i_16,
    data_arrays_1_0_reg_i_17,
    data_arrays_1_0_reg_i_18,
    data_arrays_1_0_reg_i_19,
    data_arrays_0_0_reg_i_20__0,
    data_arrays_0_0_reg_i_21__0,
    data_arrays_0_0_reg_i_22__0,
    data_arrays_0_0_reg_i_23__0,
    data_arrays_0_0_reg_i_24__0,
    data_arrays_0_0_reg_i_25__0,
    data_arrays_0_0_reg_i_26__0,
    data_arrays_0_0_reg_i_27__0,
    data_arrays_0_0_reg_i_28__0,
    tag_array_0_reg_i_8__0,
    tag_array_0_reg_i_9__0,
    tag_array_0_reg_i_10__0,
    tag_array_0_reg_i_11__0,
    tag_array_0_reg_i_12__0,
    tag_array_0_reg_i_13__0_0,
    \_T_5874_reg[1]_0 ,
    \state_reg[0] ,
    _T_5554_4_reg,
    _T_1402,
    _T_6804_0_reg,
    tile_auto_int_sync_xing_sinklzy_in_0_sync_0,
    tile_auto_int_sync_xing_sinklzy_in_0_sync_1,
    tile_auto_int_sync_xing_sinklzy_in_1_sync_0,
    q_reg,
    value_reg,
    \state_reg[0]_0 ,
    \state_reg[0]_1 ,
    \_T_1250_reg[2] ,
    \_T_5351_reg[0]_0 ,
    value_reg_0,
    _T_6059_0_reg,
    sbus_auto_coupler_from_port_named_blkdevcontroller_passthru_in_1_a_bits_address,
    resp_send_reg,
    \_T_6233_reg[5]_0 ,
    \beatsLeft_reg[1] ,
    sbus_auto_coupler_from_port_named_serialadapter_passthru_in_a_bits_address,
    \state_reg[0]_2 ,
    \_T_6233_reg[5]_1 ,
    \sendaddr_reg[11] ,
    \state_reg[0]_3 ,
    sbus_auto_coupler_from_port_named_blkdevcontroller_passthru_in_0_a_bits_address,
    _T_6418_0_reg,
    \_T_6233_reg[1]_0 ,
    \_T_5010_reg[1] ,
    maybe_full_reg_1,
    \_T_6648_reg[2] ,
    sbus_auto_coupler_to_mbus_nodelay_out_d_ready,
    \_T_558_reg[2] ,
    _T_642_0,
    _T_5577_0,
    sbus_auto_coupler_to_mbus_nodelay_out_a_bits_opcode,
    sbus_auto_coupler_from_port_named_serialadapter_passthru_in_a_bits_opcode,
    \_T_5369_reg[1] ,
    \source_reg[4] ,
    \source_reg[0] ,
    _T_920_1_reg,
    \address_reg[30] ,
    _T_920_0,
    \_T_767_reg[2]_0 ,
    count_reg_7,
    count_reg_8,
    _T_920_1,
    \address_reg[31] ,
    \address_reg[31]_0 ,
    \address_reg[31]_1 ,
    \address_reg[31]_2 ,
    io_enq_bits_param,
    io_enq_bits_source,
    io_enq_bits_data,
    \_T_1057_reg[1]_1 ,
    io_enq_bits_address,
    sys_reset_reg,
    bh_auto_out_a_ready,
    fq_reset);
  output [0:0]O;
  output mem_reg_replay_reg;
  output [8:0]ADDRARDADDR;
  output [8:0]ADDRBWRADDR;
  output [2:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_opcode;
  output [2:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_param;
  output [3:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_size;
  output [2:0]sbus_auto_coupler_to_mbus_nodelay_out_c_bits_size;
  output [0:0]DOA;
  output [3:0]\remainder_reg[107] ;
  output [3:0]\remainder_reg[111] ;
  output [3:0]\remainder_reg[115] ;
  output [0:0]\remainder_reg[115]_0 ;
  output [2:0]\remainder_reg[103] ;
  output [3:0]\remainder_reg[107]_0 ;
  output [3:0]\remainder_reg[111]_0 ;
  output [2:0]\remainder_reg[115]_1 ;
  output data_arrays_0_0_reg_i_52;
  output sbus_auto_coupler_from_tile_named_tile_fixer_in_d_ready;
  output tag_array_0_reg_i_13__0;
  output s2_valid_reg;
  output [5:0]D;
  output \_T_767_reg[2] ;
  output [1:0]\_T_5874_reg[1] ;
  output sbus_auto_coupler_from_tile_named_tile_fixer_in_a_valid;
  output [0:0]\_T_5874_reg[0] ;
  output [31:0]ram_address__T_63_data;
  output [29:0]count_reg;
  output _T_1053_reg;
  output got_e_reg;
  output got_e_reg_0;
  output [0:0]Q;
  output [0:0]\_T_5369_reg[5] ;
  output [0:0]\_T_6233_reg[5] ;
  output \_T_6215_reg[3] ;
  output \_T_6215_reg[2] ;
  output \_T_6215_reg[1] ;
  output \_T_5856_reg[0] ;
  output [0:0]\_T_5351_reg[0] ;
  output \_T_5351_reg[3] ;
  output \_T_5856_reg[3] ;
  output [0:0]DIB;
  output [0:0]\ram_opcode_reg[1] ;
  output \saved_address_reg[1] ;
  output \_T_6233_reg[0] ;
  output \saved_address_reg[1]_0 ;
  output \saved_address_reg[7] ;
  output \saved_address_reg[7]_0 ;
  output \saved_address_reg[7]_1 ;
  output \saved_address_reg[7]_2 ;
  output \saved_address_reg[7]_3 ;
  output \saved_address_reg[7]_4 ;
  output [2:0]system_bus_xbar_auto_out_3_a_bits_param;
  output [0:0]DIA;
  output [1:0]\_T_6233_reg[1] ;
  output \_T_4992_reg[2] ;
  output \_T_5874_reg[2] ;
  output \_T_6233_reg[0]_0 ;
  output _T_5195_0_reg;
  output value_1_reg;
  output \_T_4992_reg[3] ;
  output \_T_5856_reg[5] ;
  output \_T_4992_reg[7] ;
  output \_T_4992_reg[6] ;
  output \_T_4992_reg[8] ;
  output \_T_5856_reg[1] ;
  output \_T_5856_reg[2] ;
  output maybe_full_reg;
  output \_T_1057_reg[1] ;
  output \_T_1057_reg[0] ;
  output \_T_1057_reg[1]_0 ;
  output \_T_1057_reg[0]_0 ;
  output \ram_strb_reg[0] ;
  output _T_920_0_reg;
  output \ram_strb_reg[2] ;
  output \ram_strb_reg[4] ;
  output \ram_strb_reg[0]_0 ;
  output \ram_strb_reg[2]_0 ;
  output \ram_strb_reg[4]_0 ;
  output \ram_strb_reg[6] ;
  output \ram_strb_reg[6]_0 ;
  output \ram_strb_reg[1] ;
  output \ram_strb_reg[3] ;
  output \ram_strb_reg[5] ;
  output \ram_strb_reg[7] ;
  output \ram_id_reg[4] ;
  output \ram_id_reg[0] ;
  output [1:0]ram_source__T_63_data;
  output \ram_id_reg[3] ;
  output \ram_id_reg[5] ;
  output \ram_user_reg[6] ;
  output _T_940_0;
  output _T_920_3_reg;
  output maybe_full_reg_0;
  output \value_1_reg[1] ;
  output \value_1_reg[0] ;
  output _T_1670_reg;
  output _T_642_1_reg;
  output count_reg_0;
  output [0:0]count_reg_1;
  output [0:0]count_reg_2;
  output [0:0]count_reg_3;
  output [0:0]count_reg_4;
  output [0:0]count_reg_5;
  output [0:0]count_reg_6;
  output [1:0]\source_reg[1] ;
  output [7:0]ram_mask__T_63_data;
  output [63:0]ram_data__T_63_data;
  output [63:0]\ram_data_reg[63] ;
  output _GEN_61;
  output _GEN_55;
  input host_clk;
  input target_reset;
  input [2:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_opcode;
  input [3:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_size;
  input [2:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_sink;
  input sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_error;
  input tile_auto_int_sync_xing_sinklzy_in_2_sync_0;
  input [2:0]S;
  input [3:0]\remainder_reg[64] ;
  input [3:0]\remainder_reg[64]_0 ;
  input [2:0]\remainder_reg[64]_1 ;
  input [0:0]DI;
  input data_arrays_0_0_reg_i_44;
  input data_arrays_0_0_reg_i_45;
  input data_arrays_0_0_reg_i_46;
  input data_arrays_0_0_reg_i_47;
  input data_arrays_0_0_reg_i_48;
  input data_arrays_0_0_reg_i_49;
  input data_arrays_0_0_reg_i_50;
  input data_arrays_0_0_reg_i_51;
  input data_arrays_0_0_reg_i_52_0;
  input sbus_auto_coupler_from_tile_named_tile_fixer_in_b_valid;
  input sbus_auto_coupler_from_tile_named_tile_fixer_in_a_ready;
  input data_arrays_1_0_reg_i_11;
  input data_arrays_1_0_reg_i_12;
  input data_arrays_1_0_reg_i_13;
  input data_arrays_1_0_reg_i_14;
  input data_arrays_1_0_reg_i_15;
  input data_arrays_1_0_reg_i_16;
  input data_arrays_1_0_reg_i_17;
  input data_arrays_1_0_reg_i_18;
  input data_arrays_1_0_reg_i_19;
  input data_arrays_0_0_reg_i_20__0;
  input data_arrays_0_0_reg_i_21__0;
  input data_arrays_0_0_reg_i_22__0;
  input data_arrays_0_0_reg_i_23__0;
  input data_arrays_0_0_reg_i_24__0;
  input data_arrays_0_0_reg_i_25__0;
  input data_arrays_0_0_reg_i_26__0;
  input data_arrays_0_0_reg_i_27__0;
  input data_arrays_0_0_reg_i_28__0;
  input tag_array_0_reg_i_8__0;
  input tag_array_0_reg_i_9__0;
  input tag_array_0_reg_i_10__0;
  input tag_array_0_reg_i_11__0;
  input tag_array_0_reg_i_12__0;
  input tag_array_0_reg_i_13__0_0;
  input \_T_5874_reg[1]_0 ;
  input \state_reg[0] ;
  input _T_5554_4_reg;
  input _T_1402;
  input _T_6804_0_reg;
  input tile_auto_int_sync_xing_sinklzy_in_0_sync_0;
  input tile_auto_int_sync_xing_sinklzy_in_0_sync_1;
  input tile_auto_int_sync_xing_sinklzy_in_1_sync_0;
  input [0:0]q_reg;
  input value_reg;
  input \state_reg[0]_0 ;
  input \state_reg[0]_1 ;
  input \_T_1250_reg[2] ;
  input \_T_5351_reg[0]_0 ;
  input value_reg_0;
  input _T_6059_0_reg;
  input [3:0]sbus_auto_coupler_from_port_named_blkdevcontroller_passthru_in_1_a_bits_address;
  input resp_send_reg;
  input \_T_6233_reg[5]_0 ;
  input [2:0]\beatsLeft_reg[1] ;
  input [2:0]sbus_auto_coupler_from_port_named_serialadapter_passthru_in_a_bits_address;
  input \state_reg[0]_2 ;
  input \_T_6233_reg[5]_1 ;
  input [3:0]\sendaddr_reg[11] ;
  input \state_reg[0]_3 ;
  input [1:0]sbus_auto_coupler_from_port_named_blkdevcontroller_passthru_in_0_a_bits_address;
  input _T_6418_0_reg;
  input \_T_6233_reg[1]_0 ;
  input \_T_5010_reg[1] ;
  input maybe_full_reg_1;
  input \_T_6648_reg[2] ;
  input sbus_auto_coupler_to_mbus_nodelay_out_d_ready;
  input \_T_558_reg[2] ;
  input _T_642_0;
  input _T_5577_0;
  input [1:0]sbus_auto_coupler_to_mbus_nodelay_out_a_bits_opcode;
  input [0:0]sbus_auto_coupler_from_port_named_serialadapter_passthru_in_a_bits_opcode;
  input \_T_5369_reg[1] ;
  input \source_reg[4] ;
  input \source_reg[0] ;
  input _T_920_1_reg;
  input [0:0]\address_reg[30] ;
  input _T_920_0;
  input \_T_767_reg[2]_0 ;
  input count_reg_7;
  input count_reg_8;
  input _T_920_1;
  input [1:0]\address_reg[31] ;
  input [1:0]\address_reg[31]_0 ;
  input [7:0]\address_reg[31]_1 ;
  input [1:0]\address_reg[31]_2 ;
  input [1:0]io_enq_bits_param;
  input [1:0]io_enq_bits_source;
  input [63:0]io_enq_bits_data;
  input [1:0]\_T_1057_reg[1]_1 ;
  input [25:0]io_enq_bits_address;
  input sys_reset_reg;
  input bh_auto_out_a_ready;
  input fq_reset;

  wire \<const0> ;
  wire \<const1> ;
  wire [8:0]ADDRARDADDR;
  wire [8:0]ADDRBWRADDR;
  wire [5:0]D;
  wire [0:0]DI;
  wire [0:0]DIA;
  wire [0:0]DIB;
  wire [0:0]DOA;
  wire [0:0]O;
  wire [0:0]Q;
  wire \Queue/maybe_full ;
  wire \Queue/p_1_in ;
  wire \Queue/value ;
  wire \Queue/value_1 ;
  wire \Queue_3/maybe_full ;
  wire \Queue_3/value ;
  wire \Queue_3/value_1 ;
  wire [2:0]S;
  wire [63:0]_GEN_274;
  wire [126:62]_GEN_277;
  wire [31:31]_GEN_283;
  wire [25:6]_GEN_283_0;
  wire _GEN_55;
  wire _GEN_61;
  wire [6:4]_T_1005;
  wire [14:3]_T_1031;
  wire _T_1038;
  wire [5:2]_T_1050;
  wire _T_1053_reg;
  wire \_T_1057_reg[0] ;
  wire \_T_1057_reg[0]_0 ;
  wire \_T_1057_reg[1] ;
  wire \_T_1057_reg[1]_0 ;
  wire [1:0]\_T_1057_reg[1]_1 ;
  wire _T_1113;
  wire [30:12]_T_1142;
  wire _T_1156;
  wire _T_1161_1;
  wire _T_1172_1;
  wire _T_1188;
  wire [114:0]_T_1208;
  wire \_T_1250_reg[2] ;
  wire _T_1263;
  wire _T_1338;
  wire [4:0]_T_1396__T_1405_addr;
  wire [4:0]_T_1396__T_1415_addr;
  wire [2:0]_T_1396__T_2475_addr;
  wire _T_1402;
  wire [63:0]_T_1406;
  wire _T_1413;
  wire [1:0]_T_1416;
  wire _T_1488;
  wire _T_1498;
  wire _T_1573;
  wire _T_1670_reg;
  wire _T_1686;
  wire [8:0]_T_1701;
  wire _T_177;
  wire _T_179;
  wire _T_1790;
  wire _T_1821;
  wire _T_1829;
  wire _T_1844;
  wire _T_1944;
  wire _T_20810;
  wire _T_2179;
  wire _T_2181;
  wire _T_2422;
  wire _T_2425;
  wire _T_2428;
  wire _T_2431;
  wire _T_2434;
  wire _T_2437;
  wire _T_2498;
  wire _T_2499;
  wire _T_2504;
  wire _T_2507;
  wire [23:0]_T_2518;
  wire _T_2520;
  wire _T_2522;
  wire [16:16]_T_2549;
  wire _T_255;
  wire _T_258;
  wire [39:32]_T_273;
  wire [24:0]_T_2770;
  wire _T_2772;
  wire _T_2774;
  wire [1:0]_T_3585_reg__0;
  wire _T_3628;
  wire _T_384;
  wire [11:6]_T_3959;
  wire _T_407_1;
  wire _T_407_4;
  wire _T_407_6;
  wire _T_435;
  wire _T_439;
  wire _T_481;
  wire [3:3]_T_499;
  wire \_T_4992_reg[2] ;
  wire \_T_4992_reg[3] ;
  wire \_T_4992_reg[6] ;
  wire \_T_4992_reg[7] ;
  wire \_T_4992_reg[8] ;
  wire \_T_5010_reg[1] ;
  wire _T_5195_0_reg;
  wire [0:0]\_T_5351_reg[0] ;
  wire \_T_5351_reg[0]_0 ;
  wire \_T_5351_reg[3] ;
  wire \_T_5369_reg[1] ;
  wire [0:0]\_T_5369_reg[5] ;
  wire _T_5554_4_reg;
  wire _T_5577_0;
  wire \_T_558_reg[2] ;
  wire \_T_5856_reg[0] ;
  wire \_T_5856_reg[1] ;
  wire \_T_5856_reg[2] ;
  wire \_T_5856_reg[3] ;
  wire \_T_5856_reg[5] ;
  wire [0:0]\_T_5874_reg[0] ;
  wire [1:0]\_T_5874_reg[1] ;
  wire \_T_5874_reg[1]_0 ;
  wire \_T_5874_reg[2] ;
  wire _T_6059_0_reg;
  wire \_T_6215_reg[1] ;
  wire \_T_6215_reg[2] ;
  wire \_T_6215_reg[3] ;
  wire \_T_6233_reg[0] ;
  wire \_T_6233_reg[0]_0 ;
  wire [1:0]\_T_6233_reg[1] ;
  wire \_T_6233_reg[1]_0 ;
  wire [0:0]\_T_6233_reg[5] ;
  wire \_T_6233_reg[5]_0 ;
  wire \_T_6233_reg[5]_1 ;
  wire _T_628;
  wire _T_6418_0_reg;
  wire _T_642_0;
  wire _T_642_1_reg;
  wire \_T_6648_reg[2] ;
  wire _T_6804_0_reg;
  wire [63:0]_T_766;
  wire \_T_767_reg[2] ;
  wire \_T_767_reg[2]_0 ;
  wire [25:25]_T_877;
  wire [24:7]_T_889;
  wire [31:26]_T_909;
  wire _T_920_0;
  wire _T_920_0_reg;
  wire _T_920_1;
  wire _T_920_1_reg;
  wire _T_920_3_reg;
  wire _T_931;
  wire _T_940_0;
  wire _T_963;
  wire [0:0]\address_reg[30] ;
  wire [1:0]\address_reg[31] ;
  wire [1:0]\address_reg[31]_0 ;
  wire [7:0]\address_reg[31]_1 ;
  wire [1:0]\address_reg[31]_2 ;
  wire [64:64]\alu/_T_121 ;
  wire \alu/_T_217 ;
  wire \alu/_T_31 ;
  wire [5:5]\alu/shamt ;
  wire [63:15]\alu/shin ;
  wire [39:39]alu_io_adder_out;
  wire [63:1]alu_io_in1;
  wire [63:0]alu_io_in2;
  wire \arb/lastGrant ;
  wire [26:0]arb_io_out_bits_addr;
  wire [2:0]\beatsLeft_reg[1] ;
  wire bh_auto_out_a_ready;
  wire blockProbeAfterGrantCount;
  wire blockUncachedGrant;
  wire \bpu/_T_105 ;
  wire \bpu/_T_132 ;
  wire \bpu/_T_134 ;
  wire \bpu/_T_39 ;
  wire \bpu/_T_66 ;
  wire \bypass_mux_1[3]_i_7_n_0 ;
  wire \bypass_mux_1_reg[11]_i_2_n_0 ;
  wire \bypass_mux_1_reg[11]_i_2_n_1 ;
  wire \bypass_mux_1_reg[11]_i_2_n_2 ;
  wire \bypass_mux_1_reg[11]_i_2_n_3 ;
  wire \bypass_mux_1_reg[15]_i_2_n_0 ;
  wire \bypass_mux_1_reg[15]_i_2_n_1 ;
  wire \bypass_mux_1_reg[15]_i_2_n_2 ;
  wire \bypass_mux_1_reg[15]_i_2_n_3 ;
  wire \bypass_mux_1_reg[19]_i_2_n_0 ;
  wire \bypass_mux_1_reg[19]_i_2_n_1 ;
  wire \bypass_mux_1_reg[19]_i_2_n_2 ;
  wire \bypass_mux_1_reg[19]_i_2_n_3 ;
  wire \bypass_mux_1_reg[23]_i_2_n_0 ;
  wire \bypass_mux_1_reg[23]_i_2_n_1 ;
  wire \bypass_mux_1_reg[23]_i_2_n_2 ;
  wire \bypass_mux_1_reg[23]_i_2_n_3 ;
  wire \bypass_mux_1_reg[27]_i_2_n_0 ;
  wire \bypass_mux_1_reg[27]_i_2_n_1 ;
  wire \bypass_mux_1_reg[27]_i_2_n_2 ;
  wire \bypass_mux_1_reg[27]_i_2_n_3 ;
  wire \bypass_mux_1_reg[3]_i_2_n_0 ;
  wire \bypass_mux_1_reg[3]_i_2_n_1 ;
  wire \bypass_mux_1_reg[3]_i_2_n_2 ;
  wire \bypass_mux_1_reg[3]_i_2_n_3 ;
  wire \bypass_mux_1_reg[7]_i_2_n_0 ;
  wire \bypass_mux_1_reg[7]_i_2_n_1 ;
  wire \bypass_mux_1_reg[7]_i_2_n_2 ;
  wire \bypass_mux_1_reg[7]_i_2_n_3 ;
  wire \bypass_mux_2[11]_i_3_n_0 ;
  wire \bypass_mux_2[11]_i_4_n_0 ;
  wire \bypass_mux_2[11]_i_5_n_0 ;
  wire \bypass_mux_2[11]_i_6_n_0 ;
  wire \bypass_mux_2[15]_i_3_n_0 ;
  wire \bypass_mux_2[15]_i_4_n_0 ;
  wire \bypass_mux_2[15]_i_5_n_0 ;
  wire \bypass_mux_2[15]_i_6_n_0 ;
  wire \bypass_mux_2[19]_i_3_n_0 ;
  wire \bypass_mux_2[19]_i_4_n_0 ;
  wire \bypass_mux_2[19]_i_5_n_0 ;
  wire \bypass_mux_2[19]_i_6_n_0 ;
  wire \bypass_mux_2[23]_i_3_n_0 ;
  wire \bypass_mux_2[23]_i_4_n_0 ;
  wire \bypass_mux_2[23]_i_5_n_0 ;
  wire \bypass_mux_2[23]_i_6_n_0 ;
  wire \bypass_mux_2[27]_i_3_n_0 ;
  wire \bypass_mux_2[27]_i_4_n_0 ;
  wire \bypass_mux_2[27]_i_5_n_0 ;
  wire \bypass_mux_2[27]_i_6_n_0 ;
  wire \bypass_mux_2[31]_i_4_n_0 ;
  wire \bypass_mux_2[31]_i_5_n_0 ;
  wire \bypass_mux_2[31]_i_6_n_0 ;
  wire \bypass_mux_2[31]_i_7_n_0 ;
  wire \bypass_mux_2[7]_i_3_n_0 ;
  wire \bypass_mux_2[7]_i_4_n_0 ;
  wire \bypass_mux_2[7]_i_5_n_0 ;
  wire \bypass_mux_2[7]_i_6_n_0 ;
  wire \bypass_mux_2_reg[11]_i_2_n_0 ;
  wire \bypass_mux_2_reg[11]_i_2_n_1 ;
  wire \bypass_mux_2_reg[11]_i_2_n_2 ;
  wire \bypass_mux_2_reg[11]_i_2_n_3 ;
  wire \bypass_mux_2_reg[15]_i_2_n_0 ;
  wire \bypass_mux_2_reg[15]_i_2_n_1 ;
  wire \bypass_mux_2_reg[15]_i_2_n_2 ;
  wire \bypass_mux_2_reg[15]_i_2_n_3 ;
  wire \bypass_mux_2_reg[19]_i_2_n_0 ;
  wire \bypass_mux_2_reg[19]_i_2_n_1 ;
  wire \bypass_mux_2_reg[19]_i_2_n_2 ;
  wire \bypass_mux_2_reg[19]_i_2_n_3 ;
  wire \bypass_mux_2_reg[23]_i_2_n_0 ;
  wire \bypass_mux_2_reg[23]_i_2_n_1 ;
  wire \bypass_mux_2_reg[23]_i_2_n_2 ;
  wire \bypass_mux_2_reg[23]_i_2_n_3 ;
  wire \bypass_mux_2_reg[27]_i_2_n_0 ;
  wire \bypass_mux_2_reg[27]_i_2_n_1 ;
  wire \bypass_mux_2_reg[27]_i_2_n_2 ;
  wire \bypass_mux_2_reg[27]_i_2_n_3 ;
  wire \bypass_mux_2_reg[31]_i_2_n_0 ;
  wire \bypass_mux_2_reg[31]_i_2_n_1 ;
  wire \bypass_mux_2_reg[31]_i_2_n_2 ;
  wire \bypass_mux_2_reg[31]_i_2_n_3 ;
  wire \bypass_mux_2_reg[35]_i_2_n_0 ;
  wire \bypass_mux_2_reg[35]_i_2_n_1 ;
  wire \bypass_mux_2_reg[35]_i_2_n_2 ;
  wire \bypass_mux_2_reg[35]_i_2_n_3 ;
  wire \bypass_mux_2_reg[63]_i_3_n_1 ;
  wire \bypass_mux_2_reg[63]_i_3_n_2 ;
  wire \bypass_mux_2_reg[63]_i_3_n_3 ;
  wire \bypass_mux_2_reg[7]_i_2_n_0 ;
  wire \bypass_mux_2_reg[7]_i_2_n_1 ;
  wire \bypass_mux_2_reg[7]_i_2_n_2 ;
  wire \bypass_mux_2_reg[7]_i_2_n_3 ;
  wire core__100_n_0;
  wire core__101_n_0;
  wire core__102_n_0;
  wire core__103_n_0;
  wire core__104_n_0;
  wire core__105_n_0;
  wire core__106_n_0;
  wire core__107_n_0;
  wire core__108_n_0;
  wire core__109_n_0;
  wire core__10_n_0;
  wire core__110_n_0;
  wire core__111_n_0;
  wire core__112_n_0;
  wire core__113_n_0;
  wire core__114_n_0;
  wire core__115_n_0;
  wire core__116_n_0;
  wire core__117_n_0;
  wire core__118_n_0;
  wire core__119_n_0;
  wire core__11_n_0;
  wire core__120_n_0;
  wire core__121_n_0;
  wire core__122_n_0;
  wire core__123_n_0;
  wire core__124_n_0;
  wire core__125_n_0;
  wire core__126_n_0;
  wire core__127_n_0;
  wire core__128_i_14_n_0;
  wire core__128_i_14_n_1;
  wire core__128_i_14_n_2;
  wire core__128_i_14_n_3;
  wire core__128_i_19_n_0;
  wire core__128_i_19_n_1;
  wire core__128_i_19_n_2;
  wire core__128_i_19_n_3;
  wire core__128_i_28_n_0;
  wire core__128_i_28_n_1;
  wire core__128_i_28_n_2;
  wire core__128_i_28_n_3;
  wire core__128_i_33_n_0;
  wire core__128_i_33_n_1;
  wire core__128_i_33_n_2;
  wire core__128_i_33_n_3;
  wire core__128_i_3_n_1;
  wire core__128_i_3_n_2;
  wire core__128_i_3_n_3;
  wire core__128_i_46_n_0;
  wire core__128_i_46_n_1;
  wire core__128_i_46_n_2;
  wire core__128_i_46_n_3;
  wire core__128_i_4_n_0;
  wire core__128_i_4_n_1;
  wire core__128_i_4_n_2;
  wire core__128_i_4_n_3;
  wire core__128_i_6_n_0;
  wire core__128_i_6_n_1;
  wire core__128_i_6_n_2;
  wire core__128_i_6_n_3;
  wire core__128_n_0;
  wire core__129_n_0;
  wire core__12_n_0;
  wire core__130_i_4_n_0;
  wire core__130_i_4_n_1;
  wire core__130_i_4_n_2;
  wire core__130_i_4_n_3;
  wire core__130_n_0;
  wire core__131_n_0;
  wire core__132_n_0;
  wire core__133_i_3_n_0;
  wire core__133_i_3_n_1;
  wire core__133_i_3_n_2;
  wire core__133_i_3_n_3;
  wire core__133_n_0;
  wire core__134_n_0;
  wire core__135_n_0;
  wire core__136_n_0;
  wire core__137_i_3_n_0;
  wire core__137_i_3_n_1;
  wire core__137_i_3_n_2;
  wire core__137_i_3_n_3;
  wire core__137_i_3_n_4;
  wire core__137_i_3_n_5;
  wire core__137_i_3_n_6;
  wire core__137_i_3_n_7;
  wire core__137_n_0;
  wire core__138_n_0;
  wire core__139_n_0;
  wire core__13_n_0;
  wire core__140_n_0;
  wire core__141_i_3_n_0;
  wire core__141_i_3_n_1;
  wire core__141_i_3_n_2;
  wire core__141_i_3_n_3;
  wire core__141_i_3_n_4;
  wire core__141_i_3_n_5;
  wire core__141_i_3_n_6;
  wire core__141_i_3_n_7;
  wire core__141_n_0;
  wire core__142_n_0;
  wire core__143_n_0;
  wire core__144_n_0;
  wire core__145_i_4_n_0;
  wire core__145_i_4_n_1;
  wire core__145_i_4_n_2;
  wire core__145_i_4_n_3;
  wire core__145_i_4_n_4;
  wire core__145_i_4_n_5;
  wire core__145_i_4_n_6;
  wire core__145_i_4_n_7;
  wire core__145_n_0;
  wire core__146_n_0;
  wire core__147_n_0;
  wire core__148_n_0;
  wire core__149_i_4_n_0;
  wire core__149_i_4_n_1;
  wire core__149_i_4_n_2;
  wire core__149_i_4_n_3;
  wire core__149_i_4_n_4;
  wire core__149_i_4_n_5;
  wire core__149_i_4_n_6;
  wire core__149_i_4_n_7;
  wire core__149_n_0;
  wire core__14_n_0;
  wire core__150_n_0;
  wire core__151_n_0;
  wire core__152_n_0;
  wire core__153_i_4_n_0;
  wire core__153_i_4_n_1;
  wire core__153_i_4_n_2;
  wire core__153_i_4_n_3;
  wire core__153_i_4_n_4;
  wire core__153_i_4_n_5;
  wire core__153_i_4_n_6;
  wire core__153_i_4_n_7;
  wire core__153_n_0;
  wire core__154_n_0;
  wire core__155_n_0;
  wire core__156_n_0;
  wire core__157_i_3_n_1;
  wire core__157_i_3_n_2;
  wire core__157_i_3_n_3;
  wire core__157_i_3_n_4;
  wire core__157_i_3_n_5;
  wire core__157_i_3_n_6;
  wire core__157_i_3_n_7;
  wire core__157_n_0;
  wire core__158_n_0;
  wire core__159_n_0;
  wire core__15_n_0;
  wire core__160_n_0;
  wire core__161_i_1_n_0;
  wire core__161_i_1_n_1;
  wire core__161_i_1_n_2;
  wire core__161_i_1_n_3;
  wire core__161_n_0;
  wire core__162_n_0;
  wire core__163_n_0;
  wire core__164_n_0;
  wire core__165_n_0;
  wire core__166_n_0;
  wire core__167_n_0;
  wire core__168_n_0;
  wire core__169_n_0;
  wire core__16_n_0;
  wire core__170_n_0;
  wire core__171_n_0;
  wire core__172_n_0;
  wire core__173_n_0;
  wire core__174_n_0;
  wire core__175_n_0;
  wire core__176_n_0;
  wire core__177_n_0;
  wire core__178_n_0;
  wire core__179_n_0;
  wire core__17_n_0;
  wire core__180_n_0;
  wire core__181_n_0;
  wire core__182_n_0;
  wire core__183_n_0;
  wire core__184_n_0;
  wire core__185_n_0;
  wire core__186_n_0;
  wire core__187_n_0;
  wire core__188_n_0;
  wire core__189_n_0;
  wire core__18_n_0;
  wire core__190_n_0;
  wire core__191_n_0;
  wire core__192_n_0;
  wire core__193_n_0;
  wire core__194_n_0;
  wire core__195_n_0;
  wire core__196_n_0;
  wire core__197_n_0;
  wire core__198_n_0;
  wire core__199_n_0;
  wire core__19_n_0;
  wire core__200_n_0;
  wire core__201_i_1_n_0;
  wire core__201_i_1_n_1;
  wire core__201_i_1_n_2;
  wire core__201_i_1_n_3;
  wire core__201_i_2_n_0;
  wire core__201_i_3_n_0;
  wire core__201_i_4_n_0;
  wire core__201_n_0;
  wire core__202_n_0;
  wire core__203_n_0;
  wire core__204_n_0;
  wire core__205_n_0;
  wire core__206_n_0;
  wire core__207_n_0;
  wire core__208_n_0;
  wire core__209_n_0;
  wire core__20_n_0;
  wire core__210_n_0;
  wire core__211_n_0;
  wire core__212_n_0;
  wire core__213_n_0;
  wire core__214_n_0;
  wire core__215_n_0;
  wire core__216_n_0;
  wire core__217_n_0;
  wire core__218_n_0;
  wire core__219_n_0;
  wire core__21_n_0;
  wire core__220_n_0;
  wire core__221_n_0;
  wire core__222_n_0;
  wire core__223_n_0;
  wire core__224_n_0;
  wire core__225_n_0;
  wire core__226_n_0;
  wire core__227_n_0;
  wire core__228_n_0;
  wire core__229_n_0;
  wire core__22_n_0;
  wire core__230_n_0;
  wire core__231_n_0;
  wire core__232_n_0;
  wire core__233_n_0;
  wire core__234_n_0;
  wire core__235_n_0;
  wire core__236_n_0;
  wire core__237_n_0;
  wire core__238_n_0;
  wire core__239_n_0;
  wire core__23_n_0;
  wire core__240_n_0;
  wire core__241_n_0;
  wire core__242_n_0;
  wire core__243_n_0;
  wire core__244_n_0;
  wire core__245_n_0;
  wire core__246_n_0;
  wire core__247_n_0;
  wire core__248_n_0;
  wire core__249_n_0;
  wire core__24_n_0;
  wire core__250_n_0;
  wire core__251_n_0;
  wire core__252_n_0;
  wire core__253_n_0;
  wire core__254_n_0;
  wire core__255_n_0;
  wire core__256_n_0;
  wire core__257_n_0;
  wire core__258_n_0;
  wire core__259_n_0;
  wire core__25_n_0;
  wire core__260_n_0;
  wire core__261_n_0;
  wire core__262_n_0;
  wire core__263_n_0;
  wire core__264_n_0;
  wire core__265_n_0;
  wire core__266_i_11_n_0;
  wire core__266_i_11_n_1;
  wire core__266_i_11_n_2;
  wire core__266_i_11_n_3;
  wire core__266_i_16_n_0;
  wire core__266_i_16_n_1;
  wire core__266_i_16_n_2;
  wire core__266_i_16_n_3;
  wire core__266_i_1_n_3;
  wire core__266_i_21_n_0;
  wire core__266_i_21_n_1;
  wire core__266_i_21_n_2;
  wire core__266_i_21_n_3;
  wire core__266_i_3_n_0;
  wire core__266_i_3_n_1;
  wire core__266_i_3_n_2;
  wire core__266_i_3_n_3;
  wire core__266_i_4_n_0;
  wire core__266_i_6_n_0;
  wire core__266_i_6_n_1;
  wire core__266_i_6_n_2;
  wire core__266_i_6_n_3;
  wire core__266_n_0;
  wire core__267_n_0;
  wire core__268_n_0;
  wire core__269_n_0;
  wire core__26_n_0;
  wire core__270_n_0;
  wire core__271_n_0;
  wire core__272_n_0;
  wire core__273_n_0;
  wire core__274_n_0;
  wire core__275_n_0;
  wire core__276_n_0;
  wire core__277_n_0;
  wire core__278_n_0;
  wire core__279_n_0;
  wire core__27_n_0;
  wire core__280_n_0;
  wire core__281_n_0;
  wire core__282_n_0;
  wire core__283_n_0;
  wire core__284_n_0;
  wire core__285_n_0;
  wire core__286_n_0;
  wire core__287_n_0;
  wire core__288_n_0;
  wire core__289_n_0;
  wire core__28_n_0;
  wire core__290_n_0;
  wire core__291_n_0;
  wire core__292_n_0;
  wire core__293_n_0;
  wire core__294_n_0;
  wire core__295_n_0;
  wire core__296_n_0;
  wire core__297_n_0;
  wire core__298_n_0;
  wire core__299_n_0;
  wire core__29_n_0;
  wire core__300_n_0;
  wire core__301_n_0;
  wire core__302_n_0;
  wire core__303_n_0;
  wire core__304_n_0;
  wire core__305_n_0;
  wire core__306_n_0;
  wire core__307_n_0;
  wire core__308_n_0;
  wire core__309_n_0;
  wire core__30_n_0;
  wire core__310_n_0;
  wire core__311_n_0;
  wire core__312_n_0;
  wire core__313_n_0;
  wire core__314_n_0;
  wire core__315_n_0;
  wire core__316_n_0;
  wire core__317_n_0;
  wire core__318_n_0;
  wire core__319_n_0;
  wire core__31_n_0;
  wire core__320_n_0;
  wire core__321_n_0;
  wire core__322_n_0;
  wire core__323_n_0;
  wire core__324_n_0;
  wire core__325_n_0;
  wire core__326_n_0;
  wire core__327_n_0;
  wire core__328_n_0;
  wire core__329_n_0;
  wire core__32_n_0;
  wire core__330_n_0;
  wire core__331_n_0;
  wire core__332_n_0;
  wire core__333_n_0;
  wire core__334_n_0;
  wire core__335_n_0;
  wire core__336_n_0;
  wire core__337_n_0;
  wire core__338_n_0;
  wire core__339_n_0;
  wire core__33_n_0;
  wire core__340_n_0;
  wire core__341_n_0;
  wire core__342_i_10_n_0;
  wire core__342_i_12_n_0;
  wire core__342_i_13_n_0;
  wire core__342_i_14_n_0;
  wire core__342_i_15_n_0;
  wire core__342_i_20_n_0;
  wire core__342_i_21_n_0;
  wire core__342_i_22_n_0;
  wire core__342_i_23_n_0;
  wire core__342_i_4_n_0;
  wire core__342_i_5_n_0;
  wire core__342_i_6_n_0;
  wire core__342_i_8_n_0;
  wire core__342_i_9_n_0;
  wire core__342_n_0;
  wire core__343_i_2_n_0;
  wire core__343_i_3_n_0;
  wire core__343_i_4_n_0;
  wire core__343_i_5_n_0;
  wire core__343_n_0;
  wire core__344_n_0;
  wire core__345_n_0;
  wire core__346_n_0;
  wire core__347_i_2_n_0;
  wire core__347_i_3_n_0;
  wire core__347_i_4_n_0;
  wire core__347_i_5_n_0;
  wire core__347_n_0;
  wire core__348_n_0;
  wire core__349_n_0;
  wire core__34_n_0;
  wire core__350_n_0;
  wire core__351_i_2_n_0;
  wire core__351_i_3_n_0;
  wire core__351_i_4_n_0;
  wire core__351_n_0;
  wire core__352_n_0;
  wire core__353_n_0;
  wire core__354_n_0;
  wire core__355_n_0;
  wire core__356_n_0;
  wire core__357_n_0;
  wire core__358_n_0;
  wire core__359_n_0;
  wire core__35_n_0;
  wire core__360_n_0;
  wire core__361_n_0;
  wire core__362_n_0;
  wire core__363_n_0;
  wire core__364_n_0;
  wire core__365_n_0;
  wire core__366_n_0;
  wire core__367_n_0;
  wire core__368_n_0;
  wire core__369_n_0;
  wire core__36_n_0;
  wire core__370_n_0;
  wire core__371_n_0;
  wire core__372_n_0;
  wire core__373_n_0;
  wire core__374_n_0;
  wire core__375_n_0;
  wire core__376_n_0;
  wire core__377_n_0;
  wire core__378_n_0;
  wire core__379_n_0;
  wire core__37_n_0;
  wire core__380_n_0;
  wire core__381_n_0;
  wire core__382_n_0;
  wire core__383_n_0;
  wire core__384_n_0;
  wire core__385_n_0;
  wire core__386_n_0;
  wire core__387_n_0;
  wire core__388_n_0;
  wire core__389_n_0;
  wire core__38_n_0;
  wire core__390_n_0;
  wire core__391_n_0;
  wire core__392_n_0;
  wire core__393_n_0;
  wire core__394_n_0;
  wire core__395_n_0;
  wire core__396_n_0;
  wire core__397_n_0;
  wire core__398_n_0;
  wire core__399_n_0;
  wire core__39_n_0;
  wire core__400_n_0;
  wire core__401_n_0;
  wire core__402_n_0;
  wire core__403_n_0;
  wire core__404_n_0;
  wire core__405_n_0;
  wire core__406_n_0;
  wire core__407_n_0;
  wire core__408_n_0;
  wire core__409_n_0;
  wire core__40_n_0;
  wire core__410_n_0;
  wire core__411_n_0;
  wire core__412_n_0;
  wire core__413_n_0;
  wire core__414_n_0;
  wire core__415_n_0;
  wire core__416_n_0;
  wire core__417_n_0;
  wire core__418_n_0;
  wire core__419_n_0;
  wire core__41_n_0;
  wire core__420_n_0;
  wire core__421_n_0;
  wire core__422_n_0;
  wire core__423_n_0;
  wire core__424_n_0;
  wire core__425_n_0;
  wire core__426_n_0;
  wire core__427_n_0;
  wire core__428_n_0;
  wire core__429_n_0;
  wire core__42_n_0;
  wire core__430_n_0;
  wire core__431_n_0;
  wire core__432_n_0;
  wire core__433_n_0;
  wire core__434_n_0;
  wire core__435_n_0;
  wire core__436_n_0;
  wire core__437_n_0;
  wire core__438_n_0;
  wire core__439_n_0;
  wire core__43_n_0;
  wire core__440_n_0;
  wire core__441_n_0;
  wire core__442_n_0;
  wire core__443_n_0;
  wire core__444_n_0;
  wire core__445_n_0;
  wire core__446_n_0;
  wire core__447_n_0;
  wire core__448_n_0;
  wire core__449_n_0;
  wire core__44_n_0;
  wire core__450_n_0;
  wire core__451_n_0;
  wire core__452_n_0;
  wire core__453_n_0;
  wire core__454_n_0;
  wire core__455_n_0;
  wire core__456_n_0;
  wire core__457_n_0;
  wire core__458_n_0;
  wire core__459_n_0;
  wire core__45_n_0;
  wire core__460_n_0;
  wire core__461_i_10_n_0;
  wire core__461_i_10_n_1;
  wire core__461_i_10_n_2;
  wire core__461_i_10_n_3;
  wire core__461_i_5_n_0;
  wire core__461_i_5_n_1;
  wire core__461_i_5_n_2;
  wire core__461_i_5_n_3;
  wire core__461_i_7_n_0;
  wire core__461_i_7_n_1;
  wire core__461_i_7_n_2;
  wire core__461_i_7_n_3;
  wire core__461_i_9_n_0;
  wire core__461_i_9_n_1;
  wire core__461_i_9_n_2;
  wire core__461_i_9_n_3;
  wire core__462_i_10_n_2;
  wire core__462_i_10_n_3;
  wire core__462_i_11_n_2;
  wire core__462_i_11_n_3;
  wire core__462_i_12_n_2;
  wire core__462_i_12_n_3;
  wire core__462_i_3_n_2;
  wire core__462_i_3_n_3;
  wire core__462_i_4_n_2;
  wire core__462_i_4_n_3;
  wire core__462_i_5_n_2;
  wire core__462_i_5_n_3;
  wire core__462_i_6_n_2;
  wire core__462_i_6_n_3;
  wire core__462_i_7_n_2;
  wire core__462_i_7_n_3;
  wire core__462_i_8_n_2;
  wire core__462_i_8_n_3;
  wire core__462_i_9_n_2;
  wire core__462_i_9_n_3;
  wire core__46_n_0;
  wire core__47_n_0;
  wire core__48_n_0;
  wire core__49_n_0;
  wire core__4_n_0;
  wire core__501_n_0;
  wire core__502_n_0;
  wire core__503_n_0;
  wire core__504_n_0;
  wire core__505_n_0;
  wire core__506_n_0;
  wire core__507_n_0;
  wire core__508_n_0;
  wire core__509_n_0;
  wire core__50_n_0;
  wire core__510_n_0;
  wire core__51_n_0;
  wire core__52_n_0;
  wire core__53_n_0;
  wire core__54_n_0;
  wire core__550_n_0;
  wire core__551_n_0;
  wire core__552_n_0;
  wire core__553_n_0;
  wire core__554_n_0;
  wire core__555_n_0;
  wire core__556_n_0;
  wire core__557_n_0;
  wire core__558_n_0;
  wire core__55_n_0;
  wire core__56_n_0;
  wire core__57_n_0;
  wire core__58_n_0;
  wire core__598_n_0;
  wire core__59_n_0;
  wire core__5_n_0;
  wire core__60_n_0;
  wire core__61_n_0;
  wire core__62_n_0;
  wire core__638_n_0;
  wire core__639_n_0;
  wire core__63_n_0;
  wire core__640_n_0;
  wire core__641_n_0;
  wire core__642_n_0;
  wire core__643_n_0;
  wire core__644_n_0;
  wire core__645_n_0;
  wire core__646_n_0;
  wire core__647_n_0;
  wire core__648_n_0;
  wire core__649_n_0;
  wire core__64_n_0;
  wire core__650_n_0;
  wire core__651_n_0;
  wire core__652_n_0;
  wire core__653_n_0;
  wire core__654_n_0;
  wire core__655_n_0;
  wire core__656_n_0;
  wire core__657_n_0;
  wire core__658_n_0;
  wire core__659_n_0;
  wire core__65_n_0;
  wire core__660_n_0;
  wire core__661_n_0;
  wire core__662_n_0;
  wire core__663_n_0;
  wire core__664_n_0;
  wire core__665_n_0;
  wire core__666_n_0;
  wire core__667_n_0;
  wire core__668_n_0;
  wire core__669_n_0;
  wire core__66_n_0;
  wire core__670_n_0;
  wire core__671_n_0;
  wire core__672_n_0;
  wire core__673_n_0;
  wire core__674_n_0;
  wire core__675_n_0;
  wire core__676_n_0;
  wire core__677_n_0;
  wire core__678_n_0;
  wire core__679_n_0;
  wire core__67_n_0;
  wire core__680_n_0;
  wire core__681_n_0;
  wire core__682_n_0;
  wire core__683_n_0;
  wire core__684_n_0;
  wire core__685_n_0;
  wire core__686_n_0;
  wire core__687_n_0;
  wire core__688_n_0;
  wire core__68_n_0;
  wire core__691_n_0;
  wire core__692_n_0;
  wire core__695_n_0;
  wire core__697_n_0;
  wire core__698_n_0;
  wire core__699_n_0;
  wire core__69_n_0;
  wire core__6_n_0;
  wire core__702_n_0;
  wire core__704_n_0;
  wire core__705_n_0;
  wire core__706_n_0;
  wire core__708_i_12_n_0;
  wire core__708_i_16_n_0;
  wire core__708_i_16_n_1;
  wire core__708_i_16_n_2;
  wire core__708_i_16_n_3;
  wire core__708_i_21_n_0;
  wire core__708_i_21_n_1;
  wire core__708_i_21_n_2;
  wire core__708_i_21_n_3;
  wire core__708_i_30_n_0;
  wire core__708_i_30_n_1;
  wire core__708_i_30_n_2;
  wire core__708_i_30_n_3;
  wire core__708_i_35_n_0;
  wire core__708_i_35_n_1;
  wire core__708_i_35_n_2;
  wire core__708_i_35_n_3;
  wire core__708_i_48_n_0;
  wire core__708_i_48_n_1;
  wire core__708_i_48_n_2;
  wire core__708_i_48_n_3;
  wire core__708_i_5_n_1;
  wire core__708_i_5_n_2;
  wire core__708_i_5_n_3;
  wire core__708_i_6_n_0;
  wire core__708_i_6_n_1;
  wire core__708_i_6_n_2;
  wire core__708_i_6_n_3;
  wire core__708_i_8_n_0;
  wire core__708_i_8_n_1;
  wire core__708_i_8_n_2;
  wire core__708_i_8_n_3;
  wire core__708_n_0;
  wire core__709_n_0;
  wire core__70_n_0;
  wire core__710_n_0;
  wire core__714_n_0;
  wire core__715_n_0;
  wire core__716_n_0;
  wire core__717_n_0;
  wire core__71_n_0;
  wire core__72_n_0;
  wire core__73_n_0;
  wire core__74_n_0;
  wire core__75_n_0;
  wire core__76_n_0;
  wire core__77_n_0;
  wire core__78_n_0;
  wire core__79_n_0;
  wire core__7_n_0;
  wire core__80_n_0;
  wire core__81_n_0;
  wire core__82_n_0;
  wire core__83_n_0;
  wire core__84_n_0;
  wire core__85_n_0;
  wire core__86_n_0;
  wire core__87_n_0;
  wire core__88_n_0;
  wire core__89_n_0;
  wire core__8_n_0;
  wire core__90_n_0;
  wire core__91_n_0;
  wire core__92_n_0;
  wire core__93_n_0;
  wire core__94_n_0;
  wire core__95_n_0;
  wire core__96_n_0;
  wire core__97_n_0;
  wire core__98_n_0;
  wire core__99_n_0;
  wire core__9_n_0;
  wire core_n_0;
  wire core_n_1000;
  wire core_n_1001;
  wire core_n_1002;
  wire core_n_1003;
  wire core_n_1004;
  wire core_n_1005;
  wire core_n_1006;
  wire core_n_1007;
  wire core_n_1008;
  wire core_n_1009;
  wire core_n_101;
  wire core_n_1010;
  wire core_n_1011;
  wire core_n_1012;
  wire core_n_1013;
  wire core_n_1014;
  wire core_n_1015;
  wire core_n_1016;
  wire core_n_1018;
  wire core_n_1020;
  wire core_n_1028;
  wire core_n_1029;
  wire core_n_103;
  wire core_n_104;
  wire core_n_105;
  wire core_n_1069;
  wire core_n_107;
  wire core_n_1070;
  wire core_n_1071;
  wire core_n_1072;
  wire core_n_1073;
  wire core_n_1074;
  wire core_n_1075;
  wire core_n_1076;
  wire core_n_1077;
  wire core_n_1078;
  wire core_n_1079;
  wire core_n_108;
  wire core_n_1080;
  wire core_n_1081;
  wire core_n_1082;
  wire core_n_1083;
  wire core_n_1084;
  wire core_n_1085;
  wire core_n_1086;
  wire core_n_1087;
  wire core_n_1088;
  wire core_n_1089;
  wire core_n_109;
  wire core_n_1090;
  wire core_n_1091;
  wire core_n_1092;
  wire core_n_1093;
  wire core_n_1094;
  wire core_n_1095;
  wire core_n_1096;
  wire core_n_1097;
  wire core_n_1098;
  wire core_n_1099;
  wire core_n_110;
  wire core_n_1100;
  wire core_n_1102;
  wire core_n_1104;
  wire core_n_1105;
  wire core_n_1106;
  wire core_n_1107;
  wire core_n_1108;
  wire core_n_1109;
  wire core_n_111;
  wire core_n_1110;
  wire core_n_1111;
  wire core_n_1112;
  wire core_n_1113;
  wire core_n_1114;
  wire core_n_1115;
  wire core_n_1116;
  wire core_n_1117;
  wire core_n_1118;
  wire core_n_1119;
  wire core_n_112;
  wire core_n_1120;
  wire core_n_1121;
  wire core_n_1122;
  wire core_n_1128;
  wire core_n_1129;
  wire core_n_113;
  wire core_n_114;
  wire core_n_115;
  wire core_n_116;
  wire core_n_117;
  wire core_n_118;
  wire core_n_119;
  wire core_n_120;
  wire core_n_121;
  wire core_n_122;
  wire core_n_123;
  wire core_n_1238;
  wire core_n_1239;
  wire core_n_124;
  wire core_n_1240;
  wire core_n_1242;
  wire core_n_1243;
  wire core_n_1249;
  wire core_n_125;
  wire core_n_1256;
  wire core_n_1258;
  wire core_n_1259;
  wire core_n_126;
  wire core_n_1260;
  wire core_n_1261;
  wire core_n_1262;
  wire core_n_1263;
  wire core_n_1264;
  wire core_n_1265;
  wire core_n_1266;
  wire core_n_1267;
  wire core_n_1268;
  wire core_n_1269;
  wire core_n_127;
  wire core_n_1270;
  wire core_n_1271;
  wire core_n_1272;
  wire core_n_1273;
  wire core_n_1274;
  wire core_n_1275;
  wire core_n_1276;
  wire core_n_1277;
  wire core_n_128;
  wire core_n_129;
  wire core_n_130;
  wire core_n_131;
  wire core_n_1317;
  wire core_n_132;
  wire core_n_1320;
  wire core_n_1323;
  wire core_n_1329;
  wire core_n_133;
  wire core_n_1330;
  wire core_n_1331;
  wire core_n_1332;
  wire core_n_1333;
  wire core_n_1334;
  wire core_n_1335;
  wire core_n_1336;
  wire core_n_1337;
  wire core_n_1338;
  wire core_n_1339;
  wire core_n_134;
  wire core_n_1340;
  wire core_n_1341;
  wire core_n_1342;
  wire core_n_1343;
  wire core_n_1344;
  wire core_n_1345;
  wire core_n_1346;
  wire core_n_1347;
  wire core_n_1348;
  wire core_n_1349;
  wire core_n_135;
  wire core_n_1350;
  wire core_n_1354;
  wire core_n_1355;
  wire core_n_136;
  wire core_n_1360;
  wire core_n_1362;
  wire core_n_1364;
  wire core_n_1365;
  wire core_n_137;
  wire core_n_138;
  wire core_n_139;
  wire core_n_140;
  wire core_n_141;
  wire core_n_142;
  wire core_n_143;
  wire core_n_1430;
  wire core_n_1431;
  wire core_n_1432;
  wire core_n_1433;
  wire core_n_1434;
  wire core_n_1435;
  wire core_n_1436;
  wire core_n_1437;
  wire core_n_1438;
  wire core_n_1439;
  wire core_n_144;
  wire core_n_1440;
  wire core_n_1441;
  wire core_n_1442;
  wire core_n_1443;
  wire core_n_1444;
  wire core_n_1445;
  wire core_n_1446;
  wire core_n_1447;
  wire core_n_1448;
  wire core_n_1449;
  wire core_n_145;
  wire core_n_1452;
  wire core_n_1453;
  wire core_n_1454;
  wire core_n_1455;
  wire core_n_1456;
  wire core_n_1457;
  wire core_n_1458;
  wire core_n_1459;
  wire core_n_146;
  wire core_n_1460;
  wire core_n_1461;
  wire core_n_1462;
  wire core_n_1463;
  wire core_n_1464;
  wire core_n_1465;
  wire core_n_1466;
  wire core_n_1467;
  wire core_n_1468;
  wire core_n_1469;
  wire core_n_147;
  wire core_n_1470;
  wire core_n_1471;
  wire core_n_1472;
  wire core_n_1473;
  wire core_n_1474;
  wire core_n_1475;
  wire core_n_1476;
  wire core_n_1477;
  wire core_n_1478;
  wire core_n_1479;
  wire core_n_148;
  wire core_n_1480;
  wire core_n_1481;
  wire core_n_1482;
  wire core_n_1483;
  wire core_n_1484;
  wire core_n_1485;
  wire core_n_1486;
  wire core_n_1487;
  wire core_n_1488;
  wire core_n_1489;
  wire core_n_149;
  wire core_n_1490;
  wire core_n_1491;
  wire core_n_1492;
  wire core_n_1493;
  wire core_n_1494;
  wire core_n_1495;
  wire core_n_1496;
  wire core_n_1497;
  wire core_n_1498;
  wire core_n_1499;
  wire core_n_150;
  wire core_n_1500;
  wire core_n_1501;
  wire core_n_1502;
  wire core_n_1503;
  wire core_n_1504;
  wire core_n_1505;
  wire core_n_1506;
  wire core_n_1507;
  wire core_n_1508;
  wire core_n_1509;
  wire core_n_151;
  wire core_n_1510;
  wire core_n_1511;
  wire core_n_1512;
  wire core_n_1513;
  wire core_n_1514;
  wire core_n_1515;
  wire core_n_1516;
  wire core_n_1517;
  wire core_n_1518;
  wire core_n_1519;
  wire core_n_152;
  wire core_n_1520;
  wire core_n_1521;
  wire core_n_1522;
  wire core_n_1523;
  wire core_n_1524;
  wire core_n_1525;
  wire core_n_1526;
  wire core_n_1527;
  wire core_n_1528;
  wire core_n_1529;
  wire core_n_153;
  wire core_n_1530;
  wire core_n_1531;
  wire core_n_1532;
  wire core_n_1533;
  wire core_n_1534;
  wire core_n_1535;
  wire core_n_1536;
  wire core_n_1537;
  wire core_n_1538;
  wire core_n_1539;
  wire core_n_154;
  wire core_n_1540;
  wire core_n_1541;
  wire core_n_1542;
  wire core_n_1543;
  wire core_n_1544;
  wire core_n_1545;
  wire core_n_1546;
  wire core_n_1547;
  wire core_n_1548;
  wire core_n_1549;
  wire core_n_155;
  wire core_n_1550;
  wire core_n_1551;
  wire core_n_1552;
  wire core_n_1553;
  wire core_n_1554;
  wire core_n_1555;
  wire core_n_1556;
  wire core_n_1557;
  wire core_n_156;
  wire core_n_157;
  wire core_n_158;
  wire core_n_159;
  wire core_n_1591;
  wire core_n_1592;
  wire core_n_1593;
  wire core_n_1594;
  wire core_n_1595;
  wire core_n_1596;
  wire core_n_1597;
  wire core_n_1598;
  wire core_n_1599;
  wire core_n_16;
  wire core_n_160;
  wire core_n_1600;
  wire core_n_1601;
  wire core_n_1602;
  wire core_n_1603;
  wire core_n_1604;
  wire core_n_1605;
  wire core_n_1606;
  wire core_n_1607;
  wire core_n_1608;
  wire core_n_1609;
  wire core_n_161;
  wire core_n_1610;
  wire core_n_1611;
  wire core_n_1612;
  wire core_n_1613;
  wire core_n_1614;
  wire core_n_1615;
  wire core_n_162;
  wire core_n_163;
  wire core_n_164;
  wire core_n_165;
  wire core_n_166;
  wire core_n_167;
  wire core_n_168;
  wire core_n_1680;
  wire core_n_1681;
  wire core_n_1682;
  wire core_n_1683;
  wire core_n_1684;
  wire core_n_1685;
  wire core_n_1686;
  wire core_n_1687;
  wire core_n_1688;
  wire core_n_1689;
  wire core_n_169;
  wire core_n_1690;
  wire core_n_1691;
  wire core_n_1692;
  wire core_n_1693;
  wire core_n_1694;
  wire core_n_1695;
  wire core_n_1696;
  wire core_n_1697;
  wire core_n_1698;
  wire core_n_1699;
  wire core_n_1700;
  wire core_n_1701;
  wire core_n_1702;
  wire core_n_1703;
  wire core_n_1704;
  wire core_n_1705;
  wire core_n_1706;
  wire core_n_1775;
  wire core_n_1776;
  wire core_n_1777;
  wire core_n_1778;
  wire core_n_1782;
  wire core_n_1783;
  wire core_n_1784;
  wire core_n_1785;
  wire core_n_1786;
  wire core_n_1787;
  wire core_n_1788;
  wire core_n_1789;
  wire core_n_1790;
  wire core_n_1791;
  wire core_n_1792;
  wire core_n_1793;
  wire core_n_1794;
  wire core_n_1795;
  wire core_n_1796;
  wire core_n_1797;
  wire core_n_1798;
  wire core_n_1799;
  wire core_n_1800;
  wire core_n_1801;
  wire core_n_1802;
  wire core_n_1803;
  wire core_n_1804;
  wire core_n_1805;
  wire core_n_1806;
  wire core_n_1807;
  wire core_n_1808;
  wire core_n_1809;
  wire core_n_1810;
  wire core_n_1811;
  wire core_n_1812;
  wire core_n_1813;
  wire core_n_1814;
  wire core_n_1815;
  wire core_n_1816;
  wire core_n_1817;
  wire core_n_1818;
  wire core_n_1819;
  wire core_n_1820;
  wire core_n_1821;
  wire core_n_1822;
  wire core_n_1823;
  wire core_n_1824;
  wire core_n_1825;
  wire core_n_1826;
  wire core_n_1827;
  wire core_n_1828;
  wire core_n_1829;
  wire core_n_1830;
  wire core_n_1831;
  wire core_n_1832;
  wire core_n_1835;
  wire core_n_1836;
  wire core_n_1837;
  wire core_n_1838;
  wire core_n_1839;
  wire core_n_1840;
  wire core_n_1841;
  wire core_n_1842;
  wire core_n_1843;
  wire core_n_1844;
  wire core_n_1845;
  wire core_n_1846;
  wire core_n_1847;
  wire core_n_1848;
  wire core_n_1849;
  wire core_n_1850;
  wire core_n_1851;
  wire core_n_1852;
  wire core_n_1853;
  wire core_n_1854;
  wire core_n_1855;
  wire core_n_1856;
  wire core_n_1857;
  wire core_n_1858;
  wire core_n_1859;
  wire core_n_1860;
  wire core_n_1861;
  wire core_n_1862;
  wire core_n_1863;
  wire core_n_1864;
  wire core_n_1865;
  wire core_n_1866;
  wire core_n_1867;
  wire core_n_1868;
  wire core_n_1869;
  wire core_n_1870;
  wire core_n_1871;
  wire core_n_1872;
  wire core_n_1873;
  wire core_n_1874;
  wire core_n_1875;
  wire core_n_1876;
  wire core_n_1877;
  wire core_n_1878;
  wire core_n_1879;
  wire core_n_1880;
  wire core_n_1881;
  wire core_n_1882;
  wire core_n_1883;
  wire core_n_1884;
  wire core_n_1885;
  wire core_n_1886;
  wire core_n_1887;
  wire core_n_1888;
  wire core_n_1889;
  wire core_n_1890;
  wire core_n_1891;
  wire core_n_1892;
  wire core_n_1893;
  wire core_n_1894;
  wire core_n_1895;
  wire core_n_1896;
  wire core_n_1897;
  wire core_n_1898;
  wire core_n_1899;
  wire core_n_1900;
  wire core_n_1901;
  wire core_n_1902;
  wire core_n_1903;
  wire core_n_1904;
  wire core_n_1905;
  wire core_n_1906;
  wire core_n_1907;
  wire core_n_1908;
  wire core_n_1909;
  wire core_n_1910;
  wire core_n_1911;
  wire core_n_1912;
  wire core_n_1913;
  wire core_n_1914;
  wire core_n_1915;
  wire core_n_1916;
  wire core_n_1917;
  wire core_n_1918;
  wire core_n_1919;
  wire core_n_1920;
  wire core_n_1921;
  wire core_n_1922;
  wire core_n_1923;
  wire core_n_1924;
  wire core_n_1925;
  wire core_n_1926;
  wire core_n_1927;
  wire core_n_1928;
  wire core_n_1929;
  wire core_n_1930;
  wire core_n_1931;
  wire core_n_1932;
  wire core_n_1933;
  wire core_n_1934;
  wire core_n_1935;
  wire core_n_1936;
  wire core_n_1937;
  wire core_n_1938;
  wire core_n_1939;
  wire core_n_1940;
  wire core_n_1941;
  wire core_n_1942;
  wire core_n_1943;
  wire core_n_1944;
  wire core_n_1945;
  wire core_n_1946;
  wire core_n_1947;
  wire core_n_1948;
  wire core_n_1949;
  wire core_n_1950;
  wire core_n_1951;
  wire core_n_1952;
  wire core_n_1953;
  wire core_n_1954;
  wire core_n_1955;
  wire core_n_1956;
  wire core_n_1957;
  wire core_n_1958;
  wire core_n_1959;
  wire core_n_1960;
  wire core_n_1961;
  wire core_n_1962;
  wire core_n_1963;
  wire core_n_1964;
  wire core_n_1965;
  wire core_n_1966;
  wire core_n_1967;
  wire core_n_1968;
  wire core_n_1969;
  wire core_n_1970;
  wire core_n_1971;
  wire core_n_1972;
  wire core_n_1973;
  wire core_n_1974;
  wire core_n_1975;
  wire core_n_1976;
  wire core_n_1977;
  wire core_n_1978;
  wire core_n_1979;
  wire core_n_1980;
  wire core_n_1981;
  wire core_n_1982;
  wire core_n_1983;
  wire core_n_1984;
  wire core_n_1985;
  wire core_n_1986;
  wire core_n_1987;
  wire core_n_1988;
  wire core_n_1989;
  wire core_n_1990;
  wire core_n_1991;
  wire core_n_1992;
  wire core_n_1993;
  wire core_n_1994;
  wire core_n_1995;
  wire core_n_1996;
  wire core_n_1997;
  wire core_n_1998;
  wire core_n_1999;
  wire core_n_2000;
  wire core_n_2001;
  wire core_n_2002;
  wire core_n_2003;
  wire core_n_2004;
  wire core_n_2005;
  wire core_n_2006;
  wire core_n_2007;
  wire core_n_2008;
  wire core_n_2009;
  wire core_n_2010;
  wire core_n_2011;
  wire core_n_2012;
  wire core_n_2013;
  wire core_n_2014;
  wire core_n_2015;
  wire core_n_2016;
  wire core_n_2017;
  wire core_n_2018;
  wire core_n_2019;
  wire core_n_2020;
  wire core_n_2021;
  wire core_n_2022;
  wire core_n_2023;
  wire core_n_2024;
  wire core_n_2025;
  wire core_n_2026;
  wire core_n_2027;
  wire core_n_2028;
  wire core_n_2029;
  wire core_n_2030;
  wire core_n_2031;
  wire core_n_2032;
  wire core_n_2033;
  wire core_n_2034;
  wire core_n_2035;
  wire core_n_2036;
  wire core_n_2037;
  wire core_n_2038;
  wire core_n_2039;
  wire core_n_2040;
  wire core_n_2041;
  wire core_n_2042;
  wire core_n_2043;
  wire core_n_2044;
  wire core_n_2045;
  wire core_n_2046;
  wire core_n_2047;
  wire core_n_2048;
  wire core_n_2049;
  wire core_n_2050;
  wire core_n_2051;
  wire core_n_2052;
  wire core_n_2053;
  wire core_n_2054;
  wire core_n_2055;
  wire core_n_2056;
  wire core_n_2057;
  wire core_n_2058;
  wire core_n_2059;
  wire core_n_2060;
  wire core_n_2061;
  wire core_n_2062;
  wire core_n_2063;
  wire core_n_2064;
  wire core_n_2065;
  wire core_n_2066;
  wire core_n_2067;
  wire core_n_2068;
  wire core_n_2069;
  wire core_n_2070;
  wire core_n_2071;
  wire core_n_2072;
  wire core_n_2073;
  wire core_n_2074;
  wire core_n_2075;
  wire core_n_2076;
  wire core_n_2077;
  wire core_n_2078;
  wire core_n_2079;
  wire core_n_2080;
  wire core_n_2081;
  wire core_n_2082;
  wire core_n_2083;
  wire core_n_2084;
  wire core_n_2085;
  wire core_n_2086;
  wire core_n_2087;
  wire core_n_2088;
  wire core_n_2089;
  wire core_n_2090;
  wire core_n_2091;
  wire core_n_2092;
  wire core_n_2093;
  wire core_n_2094;
  wire core_n_2095;
  wire core_n_2096;
  wire core_n_2097;
  wire core_n_2098;
  wire core_n_2099;
  wire core_n_2100;
  wire core_n_2101;
  wire core_n_2102;
  wire core_n_2103;
  wire core_n_2104;
  wire core_n_2105;
  wire core_n_2106;
  wire core_n_2107;
  wire core_n_2108;
  wire core_n_2109;
  wire core_n_2110;
  wire core_n_2111;
  wire core_n_2112;
  wire core_n_2113;
  wire core_n_2114;
  wire core_n_2115;
  wire core_n_2116;
  wire core_n_2117;
  wire core_n_2118;
  wire core_n_2119;
  wire core_n_2120;
  wire core_n_2121;
  wire core_n_2122;
  wire core_n_2123;
  wire core_n_2124;
  wire core_n_2125;
  wire core_n_2126;
  wire core_n_2127;
  wire core_n_2128;
  wire core_n_2129;
  wire core_n_2130;
  wire core_n_2131;
  wire core_n_2132;
  wire core_n_2133;
  wire core_n_2134;
  wire core_n_2135;
  wire core_n_2136;
  wire core_n_2137;
  wire core_n_2138;
  wire core_n_2139;
  wire core_n_2140;
  wire core_n_2141;
  wire core_n_2142;
  wire core_n_2143;
  wire core_n_2144;
  wire core_n_2145;
  wire core_n_2146;
  wire core_n_2147;
  wire core_n_2148;
  wire core_n_2149;
  wire core_n_2150;
  wire core_n_2151;
  wire core_n_2152;
  wire core_n_2153;
  wire core_n_2154;
  wire core_n_2155;
  wire core_n_2156;
  wire core_n_2157;
  wire core_n_2158;
  wire core_n_2159;
  wire core_n_2160;
  wire core_n_2161;
  wire core_n_2162;
  wire core_n_2163;
  wire core_n_2164;
  wire core_n_2165;
  wire core_n_2166;
  wire core_n_2167;
  wire core_n_2168;
  wire core_n_2169;
  wire core_n_2170;
  wire core_n_2171;
  wire core_n_2172;
  wire core_n_2173;
  wire core_n_2174;
  wire core_n_2175;
  wire core_n_2176;
  wire core_n_2177;
  wire core_n_2178;
  wire core_n_2179;
  wire core_n_2180;
  wire core_n_2181;
  wire core_n_2182;
  wire core_n_2183;
  wire core_n_2184;
  wire core_n_2185;
  wire core_n_2186;
  wire core_n_2187;
  wire core_n_2188;
  wire core_n_2189;
  wire core_n_2190;
  wire core_n_2191;
  wire core_n_2192;
  wire core_n_2193;
  wire core_n_2194;
  wire core_n_2195;
  wire core_n_2196;
  wire core_n_2197;
  wire core_n_2198;
  wire core_n_2199;
  wire core_n_2200;
  wire core_n_2201;
  wire core_n_2203;
  wire core_n_2204;
  wire core_n_2205;
  wire core_n_2206;
  wire core_n_2207;
  wire core_n_2208;
  wire core_n_2209;
  wire core_n_2210;
  wire core_n_2211;
  wire core_n_2212;
  wire core_n_2213;
  wire core_n_2214;
  wire core_n_2215;
  wire core_n_2216;
  wire core_n_2217;
  wire core_n_2218;
  wire core_n_2219;
  wire core_n_2220;
  wire core_n_2221;
  wire core_n_2222;
  wire core_n_2223;
  wire core_n_2224;
  wire core_n_2225;
  wire core_n_2226;
  wire core_n_2227;
  wire core_n_2228;
  wire core_n_2229;
  wire core_n_2230;
  wire core_n_2231;
  wire core_n_2232;
  wire core_n_2233;
  wire core_n_2234;
  wire core_n_2240;
  wire core_n_2241;
  wire core_n_2242;
  wire core_n_2243;
  wire core_n_2244;
  wire core_n_2245;
  wire core_n_2246;
  wire core_n_2247;
  wire core_n_2248;
  wire core_n_2249;
  wire core_n_2250;
  wire core_n_2251;
  wire core_n_2252;
  wire core_n_2253;
  wire core_n_2254;
  wire core_n_2255;
  wire core_n_2256;
  wire core_n_2257;
  wire core_n_2259;
  wire core_n_2260;
  wire core_n_2261;
  wire core_n_2262;
  wire core_n_2263;
  wire core_n_2264;
  wire core_n_2265;
  wire core_n_2266;
  wire core_n_2267;
  wire core_n_2268;
  wire core_n_2269;
  wire core_n_2270;
  wire core_n_2271;
  wire core_n_2272;
  wire core_n_2273;
  wire core_n_2274;
  wire core_n_2275;
  wire core_n_2276;
  wire core_n_2277;
  wire core_n_2278;
  wire core_n_2279;
  wire core_n_2280;
  wire core_n_2281;
  wire core_n_2282;
  wire core_n_2283;
  wire core_n_2284;
  wire core_n_2285;
  wire core_n_2286;
  wire core_n_2287;
  wire core_n_2288;
  wire core_n_2289;
  wire core_n_2290;
  wire core_n_2291;
  wire core_n_2292;
  wire core_n_2293;
  wire core_n_2294;
  wire core_n_2295;
  wire core_n_2296;
  wire core_n_2297;
  wire core_n_2298;
  wire core_n_2299;
  wire core_n_2300;
  wire core_n_2301;
  wire core_n_2302;
  wire core_n_2303;
  wire core_n_2304;
  wire core_n_2305;
  wire core_n_2306;
  wire core_n_2307;
  wire core_n_2308;
  wire core_n_2309;
  wire core_n_2310;
  wire core_n_2311;
  wire core_n_2312;
  wire core_n_2313;
  wire core_n_2314;
  wire core_n_2315;
  wire core_n_2316;
  wire core_n_2317;
  wire core_n_2318;
  wire core_n_2319;
  wire core_n_2320;
  wire core_n_2321;
  wire core_n_2322;
  wire core_n_2323;
  wire core_n_2324;
  wire core_n_2325;
  wire core_n_2326;
  wire core_n_2327;
  wire core_n_2328;
  wire core_n_2329;
  wire core_n_237;
  wire core_n_238;
  wire core_n_265;
  wire core_n_266;
  wire core_n_267;
  wire core_n_268;
  wire core_n_269;
  wire core_n_270;
  wire core_n_271;
  wire core_n_272;
  wire core_n_273;
  wire core_n_274;
  wire core_n_275;
  wire core_n_276;
  wire core_n_277;
  wire core_n_278;
  wire core_n_279;
  wire core_n_28;
  wire core_n_280;
  wire core_n_281;
  wire core_n_282;
  wire core_n_283;
  wire core_n_284;
  wire core_n_285;
  wire core_n_286;
  wire core_n_287;
  wire core_n_288;
  wire core_n_289;
  wire core_n_30;
  wire core_n_310;
  wire core_n_32;
  wire core_n_323;
  wire core_n_324;
  wire core_n_325;
  wire core_n_327;
  wire core_n_328;
  wire core_n_329;
  wire core_n_330;
  wire core_n_331;
  wire core_n_332;
  wire core_n_333;
  wire core_n_334;
  wire core_n_335;
  wire core_n_336;
  wire core_n_337;
  wire core_n_338;
  wire core_n_339;
  wire core_n_340;
  wire core_n_341;
  wire core_n_342;
  wire core_n_343;
  wire core_n_344;
  wire core_n_345;
  wire core_n_346;
  wire core_n_347;
  wire core_n_348;
  wire core_n_349;
  wire core_n_350;
  wire core_n_351;
  wire core_n_352;
  wire core_n_353;
  wire core_n_354;
  wire core_n_356;
  wire core_n_357;
  wire core_n_358;
  wire core_n_359;
  wire core_n_360;
  wire core_n_361;
  wire core_n_362;
  wire core_n_363;
  wire core_n_364;
  wire core_n_365;
  wire core_n_366;
  wire core_n_367;
  wire core_n_368;
  wire core_n_369;
  wire core_n_370;
  wire core_n_371;
  wire core_n_372;
  wire core_n_373;
  wire core_n_374;
  wire core_n_375;
  wire core_n_387;
  wire core_n_391;
  wire core_n_392;
  wire core_n_393;
  wire core_n_423;
  wire core_n_424;
  wire core_n_425;
  wire core_n_426;
  wire core_n_459;
  wire core_n_518;
  wire core_n_519;
  wire core_n_520;
  wire core_n_551;
  wire core_n_639;
  wire core_n_640;
  wire core_n_641;
  wire core_n_642;
  wire core_n_643;
  wire core_n_644;
  wire core_n_645;
  wire core_n_646;
  wire core_n_647;
  wire core_n_649;
  wire core_n_651;
  wire core_n_652;
  wire core_n_68;
  wire core_n_680;
  wire core_n_682;
  wire core_n_685;
  wire core_n_686;
  wire core_n_687;
  wire core_n_69;
  wire core_n_692;
  wire core_n_693;
  wire core_n_694;
  wire core_n_695;
  wire core_n_70;
  wire core_n_700;
  wire core_n_701;
  wire core_n_702;
  wire core_n_703;
  wire core_n_708;
  wire core_n_709;
  wire core_n_710;
  wire core_n_711;
  wire core_n_712;
  wire core_n_713;
  wire core_n_714;
  wire core_n_715;
  wire core_n_721;
  wire core_n_722;
  wire core_n_723;
  wire core_n_724;
  wire core_n_730;
  wire core_n_731;
  wire core_n_732;
  wire core_n_733;
  wire core_n_736;
  wire core_n_737;
  wire core_n_738;
  wire core_n_739;
  wire core_n_745;
  wire core_n_746;
  wire core_n_747;
  wire core_n_748;
  wire core_n_749;
  wire core_n_752;
  wire core_n_753;
  wire core_n_754;
  wire core_n_755;
  wire core_n_756;
  wire core_n_757;
  wire core_n_758;
  wire core_n_759;
  wire core_n_760;
  wire core_n_761;
  wire core_n_762;
  wire core_n_763;
  wire core_n_764;
  wire core_n_765;
  wire core_n_766;
  wire core_n_767;
  wire core_n_768;
  wire core_n_769;
  wire core_n_770;
  wire core_n_771;
  wire core_n_772;
  wire core_n_773;
  wire core_n_774;
  wire core_n_775;
  wire core_n_776;
  wire core_n_777;
  wire core_n_778;
  wire core_n_779;
  wire core_n_780;
  wire core_n_781;
  wire core_n_782;
  wire core_n_783;
  wire core_n_784;
  wire core_n_785;
  wire core_n_786;
  wire core_n_787;
  wire core_n_788;
  wire core_n_789;
  wire core_n_790;
  wire core_n_791;
  wire core_n_792;
  wire core_n_793;
  wire core_n_794;
  wire core_n_795;
  wire core_n_796;
  wire core_n_797;
  wire core_n_798;
  wire core_n_799;
  wire core_n_800;
  wire core_n_801;
  wire core_n_802;
  wire core_n_803;
  wire core_n_804;
  wire core_n_805;
  wire core_n_806;
  wire core_n_807;
  wire core_n_808;
  wire core_n_809;
  wire core_n_811;
  wire core_n_812;
  wire core_n_813;
  wire core_n_814;
  wire core_n_815;
  wire core_n_816;
  wire core_n_817;
  wire core_n_818;
  wire core_n_819;
  wire core_n_82;
  wire core_n_820;
  wire core_n_821;
  wire core_n_822;
  wire core_n_823;
  wire core_n_824;
  wire core_n_825;
  wire core_n_826;
  wire core_n_827;
  wire core_n_828;
  wire core_n_829;
  wire core_n_830;
  wire core_n_831;
  wire core_n_832;
  wire core_n_833;
  wire core_n_834;
  wire core_n_835;
  wire core_n_836;
  wire core_n_837;
  wire core_n_838;
  wire core_n_839;
  wire core_n_840;
  wire core_n_841;
  wire core_n_842;
  wire core_n_843;
  wire core_n_844;
  wire core_n_845;
  wire core_n_846;
  wire core_n_847;
  wire core_n_848;
  wire core_n_849;
  wire core_n_85;
  wire core_n_850;
  wire core_n_851;
  wire core_n_852;
  wire core_n_853;
  wire core_n_854;
  wire core_n_855;
  wire core_n_856;
  wire core_n_857;
  wire core_n_858;
  wire core_n_859;
  wire core_n_86;
  wire core_n_860;
  wire core_n_861;
  wire core_n_862;
  wire core_n_863;
  wire core_n_864;
  wire core_n_865;
  wire core_n_866;
  wire core_n_867;
  wire core_n_868;
  wire core_n_869;
  wire core_n_870;
  wire core_n_871;
  wire core_n_872;
  wire core_n_873;
  wire core_n_874;
  wire core_n_875;
  wire core_n_876;
  wire core_n_877;
  wire core_n_878;
  wire core_n_879;
  wire core_n_880;
  wire core_n_881;
  wire core_n_882;
  wire core_n_883;
  wire core_n_884;
  wire core_n_885;
  wire core_n_886;
  wire core_n_887;
  wire core_n_888;
  wire core_n_889;
  wire core_n_890;
  wire core_n_891;
  wire core_n_892;
  wire core_n_894;
  wire core_n_895;
  wire core_n_896;
  wire core_n_897;
  wire core_n_901;
  wire core_n_902;
  wire core_n_904;
  wire core_n_906;
  wire core_n_907;
  wire core_n_908;
  wire core_n_909;
  wire core_n_91;
  wire core_n_910;
  wire core_n_912;
  wire core_n_913;
  wire core_n_914;
  wire core_n_92;
  wire core_n_93;
  wire core_n_940;
  wire core_n_941;
  wire core_n_942;
  wire core_n_943;
  wire core_n_944;
  wire core_n_945;
  wire core_n_946;
  wire core_n_947;
  wire core_n_948;
  wire core_n_949;
  wire core_n_95;
  wire core_n_950;
  wire core_n_951;
  wire core_n_952;
  wire core_n_953;
  wire core_n_954;
  wire core_n_955;
  wire core_n_956;
  wire core_n_957;
  wire core_n_958;
  wire core_n_959;
  wire core_n_962;
  wire core_n_963;
  wire core_n_964;
  wire core_n_965;
  wire core_n_966;
  wire core_n_968;
  wire core_n_969;
  wire core_n_970;
  wire core_n_971;
  wire core_n_972;
  wire core_n_973;
  wire core_n_974;
  wire core_n_975;
  wire core_n_976;
  wire core_n_977;
  wire core_n_98;
  wire core_n_99;
  wire core_n_992;
  wire core_n_994;
  wire core_n_995;
  wire core_n_996;
  wire core_n_997;
  wire core_n_999;
  wire core_rep__0_n_0;
  wire core_rep__10_n_0;
  wire core_rep__11_n_0;
  wire core_rep__12_n_0;
  wire core_rep__13_n_0;
  wire core_rep__14_n_0;
  wire core_rep__15_n_0;
  wire core_rep__16_n_0;
  wire core_rep__17_n_0;
  wire core_rep__18_n_0;
  wire core_rep__19_n_0;
  wire core_rep__1_n_0;
  wire core_rep__20_n_0;
  wire core_rep__21_n_0;
  wire core_rep__22_n_0;
  wire core_rep__23_n_0;
  wire core_rep__24_n_0;
  wire core_rep__25_n_0;
  wire core_rep__26_n_0;
  wire core_rep__27_n_0;
  wire core_rep__28_n_0;
  wire core_rep__29_n_0;
  wire core_rep__2_n_0;
  wire core_rep__30_n_0;
  wire core_rep__31_n_0;
  wire core_rep__32_n_0;
  wire core_rep__33_n_0;
  wire core_rep__34_n_0;
  wire core_rep__35_n_0;
  wire core_rep__36_n_0;
  wire core_rep__3_n_0;
  wire core_rep__4_n_0;
  wire core_rep__5_n_0;
  wire core_rep__6_n_0;
  wire core_rep__7_n_0;
  wire core_rep__8_n_0;
  wire core_rep__9_n_0;
  wire core_rep_n_0;
  wire [29:0]count_reg;
  wire count_reg_0;
  wire [0:0]count_reg_1;
  wire [0:0]count_reg_2;
  wire [0:0]count_reg_3;
  wire [0:0]count_reg_4;
  wire [0:0]count_reg_5;
  wire [0:0]count_reg_6;
  wire count_reg_7;
  wire count_reg_8;
  wire [39:1]\csr/_GEN_350 ;
  wire [39:1]\csr/_GEN_364 ;
  wire [39:1]\csr/_GEN_369 ;
  wire [6:6]\csr/_T_286__0 ;
  wire [39:5]\csr/_T_4899 ;
  wire [63:0]\csr/_T_5044 ;
  wire \csr/_T_5074 ;
  wire [39:0]\csr/p_1_in ;
  wire \csr/reg_dcsr_prv ;
  wire \csr/reg_dcsr_step ;
  wire \csr/reg_mstatus_mie ;
  wire [4:4]\csr/reg_mtvec ;
  wire \csr/reg_singleStepped ;
  wire [4:4]\csr/reg_stvec ;
  wire [38:0]csr_io_bp_0_address;
  wire csr_io_bp_0_control_action;
  wire csr_io_bp_0_control_m;
  wire csr_io_bp_0_control_s;
  wire [0:0]csr_io_bp_0_control_tmatch;
  wire csr_io_bp_0_control_u;
  wire [11:0]csr_io_rw_addr;
  wire csr_io_status_debug;
  wire [12:2]csr_io_status_isa;
  wire [39:39]csr_io_tval;
  wire [11:6]dataArb_io_in_1_bits_addr;
  wire dataArb_io_in_1_valid;
  wire dataArb_io_in_2_valid;
  wire data_arrays_0_0_reg_i_20__0;
  wire data_arrays_0_0_reg_i_21__0;
  wire data_arrays_0_0_reg_i_22__0;
  wire data_arrays_0_0_reg_i_23__0;
  wire data_arrays_0_0_reg_i_24__0;
  wire data_arrays_0_0_reg_i_25__0;
  wire data_arrays_0_0_reg_i_26__0;
  wire data_arrays_0_0_reg_i_27__0;
  wire data_arrays_0_0_reg_i_28__0;
  wire data_arrays_0_0_reg_i_44;
  wire data_arrays_0_0_reg_i_45;
  wire data_arrays_0_0_reg_i_46;
  wire data_arrays_0_0_reg_i_47;
  wire data_arrays_0_0_reg_i_48;
  wire data_arrays_0_0_reg_i_49;
  wire data_arrays_0_0_reg_i_50;
  wire data_arrays_0_0_reg_i_51;
  wire data_arrays_0_0_reg_i_52;
  wire data_arrays_0_0_reg_i_52_0;
  wire data_arrays_1_0_reg_i_11;
  wire data_arrays_1_0_reg_i_12;
  wire data_arrays_1_0_reg_i_13;
  wire data_arrays_1_0_reg_i_14;
  wire data_arrays_1_0_reg_i_15;
  wire data_arrays_1_0_reg_i_16;
  wire data_arrays_1_0_reg_i_17;
  wire data_arrays_1_0_reg_i_18;
  wire data_arrays_1_0_reg_i_19;
  wire [11:3]dcacheArb_io_requestor_0_req_bits_addr;
  wire dcacheArb_io_requestor_0_req_ready;
  wire dcacheArb_io_requestor_0_s1_kill;
  wire dcacheArb_io_requestor_1_ordered;
  wire dcacheArb_io_requestor_1_replay_next;
  wire [38:0]dcacheArb_io_requestor_1_req_bits_addr;
  wire [4:0]dcacheArb_io_requestor_1_req_bits_cmd;
  wire [5:1]dcacheArb_io_requestor_1_req_bits_tag;
  wire [2:0]dcacheArb_io_requestor_1_req_bits_typ;
  wire dcacheArb_io_requestor_1_req_ready;
  wire dcacheArb_io_requestor_1_req_valid;
  wire [63:0]dcacheArb_io_requestor_1_resp_bits_data;
  wire [63:0]dcacheArb_io_requestor_1_resp_bits_data_word_bypass;
  wire dcacheArb_io_requestor_1_resp_bits_replay;
  wire [5:1]dcacheArb_io_requestor_1_resp_bits_tag;
  wire dcacheArb_io_requestor_1_resp_valid;
  wire [63:0]dcacheArb_io_requestor_1_s1_data_data;
  wire dcacheArb_io_requestor_1_s1_kill;
  wire dcacheArb_io_requestor_1_s2_nack;
  wire dcacheArb_io_requestor_1_s2_xcpt_ae_ld;
  wire dcacheArb_io_requestor_1_s2_xcpt_ma_ld;
  wire dcacheArb_io_requestor_1_s2_xcpt_ma_st;
  wire dcacheArb_io_requestor_1_s2_xcpt_pf_ld;
  wire dcacheArb_io_requestor_1_s2_xcpt_pf_st;
  wire dcache_io_cpu_invalidate_lr;
  wire [31:3]dcache_io_cpu_req_bits_addr;
  wire [26:0]dcache_io_ptw_req_bits_addr;
  wire dcache_io_ptw_resp_bits_ae;
  wire dcache_io_ptw_resp_bits_homogeneous;
  wire [1:0]dcache_io_ptw_resp_bits_level;
  wire dcache_io_ptw_resp_bits_pte_g;
  wire [19:0]dcache_io_ptw_resp_bits_pte_ppn;
  wire dcache_io_ptw_resp_bits_pte_u;
  wire dcache_io_ptw_resp_bits_pte_v;
  wire dcache_io_ptw_resp_valid;
  wire [1:0]dcache_io_ptw_status_dprv;
  wire dcache_io_ptw_status_mxr;
  wire dcache_io_ptw_status_sum;
  wire dcache_n_0;
  wire dcache_n_1;
  wire dcache_n_133;
  wire dcache_n_134;
  wire dcache_n_136;
  wire dcache_n_137;
  wire dcache_n_138;
  wire dcache_n_139;
  wire dcache_n_140;
  wire dcache_n_141;
  wire dcache_n_142;
  wire dcache_n_143;
  wire dcache_n_144;
  wire dcache_n_145;
  wire dcache_n_146;
  wire dcache_n_147;
  wire dcache_n_148;
  wire dcache_n_149;
  wire dcache_n_150;
  wire dcache_n_151;
  wire dcache_n_152;
  wire dcache_n_153;
  wire dcache_n_154;
  wire dcache_n_155;
  wire dcache_n_156;
  wire dcache_n_157;
  wire dcache_n_158;
  wire dcache_n_159;
  wire dcache_n_161;
  wire dcache_n_17;
  wire dcache_n_18;
  wire dcache_n_19;
  wire dcache_n_2;
  wire dcache_n_20;
  wire dcache_n_209;
  wire dcache_n_21;
  wire dcache_n_210;
  wire dcache_n_212;
  wire dcache_n_213;
  wire dcache_n_22;
  wire dcache_n_23;
  wire dcache_n_24;
  wire dcache_n_25;
  wire dcache_n_26;
  wire dcache_n_27;
  wire dcache_n_28;
  wire dcache_n_29;
  wire dcache_n_3;
  wire dcache_n_30;
  wire dcache_n_31;
  wire dcache_n_32;
  wire dcache_n_33;
  wire dcache_n_34;
  wire dcache_n_342;
  wire dcache_n_343;
  wire dcache_n_346;
  wire dcache_n_35;
  wire dcache_n_36;
  wire dcache_n_367;
  wire dcache_n_368;
  wire dcache_n_369;
  wire dcache_n_37;
  wire dcache_n_370;
  wire dcache_n_371;
  wire dcache_n_372;
  wire dcache_n_373;
  wire dcache_n_374;
  wire dcache_n_375;
  wire dcache_n_376;
  wire dcache_n_377;
  wire dcache_n_378;
  wire dcache_n_379;
  wire dcache_n_38;
  wire dcache_n_380;
  wire dcache_n_381;
  wire dcache_n_382;
  wire dcache_n_383;
  wire dcache_n_384;
  wire dcache_n_385;
  wire dcache_n_386;
  wire dcache_n_387;
  wire dcache_n_388;
  wire dcache_n_39;
  wire dcache_n_4;
  wire dcache_n_40;
  wire dcache_n_41;
  wire dcache_n_415;
  wire dcache_n_416;
  wire dcache_n_417;
  wire dcache_n_418;
  wire dcache_n_42;
  wire dcache_n_423;
  wire dcache_n_429;
  wire dcache_n_43;
  wire dcache_n_431;
  wire dcache_n_432;
  wire dcache_n_433;
  wire dcache_n_435;
  wire dcache_n_436;
  wire dcache_n_438;
  wire dcache_n_439;
  wire dcache_n_44;
  wire dcache_n_440;
  wire dcache_n_441;
  wire dcache_n_442;
  wire dcache_n_443;
  wire dcache_n_448;
  wire dcache_n_45;
  wire dcache_n_453;
  wire dcache_n_454;
  wire dcache_n_455;
  wire dcache_n_456;
  wire dcache_n_46;
  wire dcache_n_47;
  wire dcache_n_48;
  wire dcache_n_49;
  wire dcache_n_5;
  wire dcache_n_50;
  wire dcache_n_51;
  wire dcache_n_52;
  wire dcache_n_53;
  wire dcache_n_54;
  wire dcache_n_541;
  wire dcache_n_542;
  wire dcache_n_543;
  wire dcache_n_544;
  wire dcache_n_55;
  wire dcache_n_550;
  wire dcache_n_551;
  wire dcache_n_552;
  wire dcache_n_553;
  wire dcache_n_554;
  wire dcache_n_555;
  wire dcache_n_556;
  wire dcache_n_557;
  wire dcache_n_558;
  wire dcache_n_559;
  wire dcache_n_56;
  wire dcache_n_560;
  wire dcache_n_561;
  wire dcache_n_562;
  wire dcache_n_563;
  wire dcache_n_564;
  wire dcache_n_565;
  wire dcache_n_566;
  wire dcache_n_567;
  wire dcache_n_569;
  wire dcache_n_57;
  wire dcache_n_570;
  wire dcache_n_571;
  wire dcache_n_572;
  wire dcache_n_573;
  wire dcache_n_574;
  wire dcache_n_575;
  wire dcache_n_576;
  wire dcache_n_578;
  wire dcache_n_58;
  wire dcache_n_580;
  wire dcache_n_582;
  wire dcache_n_583;
  wire dcache_n_584;
  wire dcache_n_585;
  wire dcache_n_59;
  wire dcache_n_6;
  wire dcache_n_60;
  wire dcache_n_61;
  wire dcache_n_610;
  wire dcache_n_611;
  wire dcache_n_612;
  wire dcache_n_613;
  wire dcache_n_614;
  wire dcache_n_615;
  wire dcache_n_616;
  wire dcache_n_617;
  wire dcache_n_618;
  wire dcache_n_619;
  wire dcache_n_62;
  wire dcache_n_620;
  wire dcache_n_621;
  wire dcache_n_622;
  wire dcache_n_623;
  wire dcache_n_624;
  wire dcache_n_625;
  wire dcache_n_626;
  wire dcache_n_627;
  wire dcache_n_628;
  wire dcache_n_629;
  wire dcache_n_63;
  wire dcache_n_630;
  wire dcache_n_631;
  wire dcache_n_632;
  wire dcache_n_633;
  wire dcache_n_634;
  wire dcache_n_635;
  wire dcache_n_636;
  wire dcache_n_637;
  wire dcache_n_638;
  wire dcache_n_639;
  wire dcache_n_64;
  wire dcache_n_640;
  wire dcache_n_641;
  wire dcache_n_642;
  wire dcache_n_643;
  wire dcache_n_65;
  wire dcache_n_66;
  wire dcache_n_67;
  wire dcache_n_68;
  wire dcache_n_69;
  wire dcache_n_7;
  wire dcache_n_70;
  wire dcache_n_71;
  wire dcache_n_72;
  wire dcache_n_75;
  wire dcache_n_89;
  wire dcache_n_90;
  wire [1:0]\div/_GEN_35 ;
  wire [63:0]\div/_GEN_36 ;
  wire \div/_T_103 ;
  wire [61:61]\div/_T_122 ;
  wire [0:0]\div/_T_216 ;
  wire [9:9]\div/_T_94 ;
  wire [9:9]\div/p_1_in ;
  wire [29:10]div_io_resp_bits_data;
  wire [4:0]div_io_resp_bits_tag;
  wire [3:3]ex_ctrl_alu_fn;
  wire ex_ctrl_div;
  wire ex_ctrl_fence_i;
  wire ex_ctrl_jalr;
  wire [1:0]ex_ctrl_sel_alu2;
  wire [2:0]ex_ctrl_sel_imm;
  wire ex_ctrl_wxd;
  wire ex_reg_flush_pipe;
  wire [31:31]ex_reg_pc;
  wire [1:0]ex_reg_rs_lsb_1;
  wire ex_reg_rs_msb_0;
  wire ex_reg_valid;
  wire ex_reg_xcpt;
  wire ex_reg_xcpt_interrupt;
  wire ex_sfence;
  wire [38:38]\fq/elts_0_pc ;
  wire [2:2]fq_io_mask;
  wire fq_reset;
  wire [39:2]frontend_io_cpu_req_bits_pc;
  wire frontend_io_cpu_req_bits_speculative;
  wire [30:3]frontend_io_cpu_resp_bits_data;
  wire [39:1]frontend_io_cpu_resp_bits_pc;
  wire frontend_io_cpu_resp_bits_replay;
  wire frontend_io_cpu_resp_bits_xcpt_ae_inst;
  wire frontend_io_cpu_resp_bits_xcpt_pf_inst;
  wire frontend_io_cpu_resp_valid;
  wire frontend_io_cpu_sfence_bits_rs1;
  wire frontend_io_cpu_sfence_valid;
  wire [29:0]frontend_io_ptw_pmp_0_addr;
  wire [29:0]frontend_io_ptw_pmp_1_addr;
  wire [1:0]frontend_io_ptw_pmp_1_cfg_a;
  wire frontend_io_ptw_pmp_1_cfg_w;
  wire [29:11]frontend_io_ptw_pmp_1_mask;
  wire [29:0]frontend_io_ptw_pmp_2_addr;
  wire [1:0]frontend_io_ptw_pmp_2_cfg_a;
  wire [29:11]frontend_io_ptw_pmp_2_mask;
  wire [29:0]frontend_io_ptw_pmp_3_addr;
  wire [29:0]frontend_io_ptw_pmp_4_addr;
  wire [1:1]frontend_io_ptw_pmp_4_cfg_a;
  wire [29:11]frontend_io_ptw_pmp_4_mask;
  wire [29:0]frontend_io_ptw_pmp_5_addr;
  wire [1:1]frontend_io_ptw_pmp_5_cfg_a;
  wire [29:11]frontend_io_ptw_pmp_5_mask;
  wire [29:0]frontend_io_ptw_pmp_6_addr;
  wire [1:0]frontend_io_ptw_pmp_6_cfg_a;
  wire [29:11]frontend_io_ptw_pmp_6_mask;
  wire [29:0]frontend_io_ptw_pmp_7_addr;
  wire [1:0]frontend_io_ptw_pmp_7_cfg_a;
  wire [29:11]frontend_io_ptw_pmp_7_mask;
  wire [3:3]frontend_io_ptw_ptbr_mode;
  wire frontend_io_ptw_req_ready;
  wire [1:0]frontend_io_ptw_status_prv;
  wire frontend_n_114;
  wire frontend_n_115;
  wire frontend_n_116;
  wire frontend_n_117;
  wire frontend_n_118;
  wire frontend_n_119;
  wire frontend_n_120;
  wire frontend_n_121;
  wire frontend_n_125;
  wire frontend_n_126;
  wire frontend_n_127;
  wire frontend_n_128;
  wire frontend_n_129;
  wire frontend_n_130;
  wire frontend_n_131;
  wire frontend_n_132;
  wire frontend_n_133;
  wire frontend_n_134;
  wire frontend_n_136;
  wire frontend_n_137;
  wire frontend_n_138;
  wire frontend_n_139;
  wire frontend_n_140;
  wire frontend_n_141;
  wire frontend_n_142;
  wire frontend_n_143;
  wire frontend_n_144;
  wire frontend_n_145;
  wire frontend_n_146;
  wire frontend_n_147;
  wire frontend_n_148;
  wire frontend_n_149;
  wire frontend_n_150;
  wire frontend_n_151;
  wire frontend_n_152;
  wire frontend_n_169;
  wire frontend_n_170;
  wire frontend_n_222;
  wire frontend_n_223;
  wire frontend_n_224;
  wire frontend_n_225;
  wire frontend_n_226;
  wire frontend_n_230;
  wire frontend_n_231;
  wire frontend_n_232;
  wire frontend_n_239;
  wire frontend_n_240;
  wire frontend_n_241;
  wire frontend_n_243;
  wire frontend_n_244;
  wire frontend_n_245;
  wire frontend_n_265;
  wire frontend_n_267;
  wire frontend_n_268;
  wire frontend_n_269;
  wire frontend_n_285;
  wire frontend_n_293;
  wire frontend_n_294;
  wire frontend_n_300;
  wire frontend_n_304;
  wire frontend_n_312;
  wire frontend_n_318;
  wire frontend_n_320;
  wire frontend_n_351;
  wire frontend_n_352;
  wire frontend_n_353;
  wire frontend_n_354;
  wire frontend_n_355;
  wire frontend_n_356;
  wire frontend_n_358;
  wire frontend_n_359;
  wire frontend_n_360;
  wire frontend_n_361;
  wire frontend_n_362;
  wire frontend_n_364;
  wire frontend_n_365;
  wire frontend_n_366;
  wire frontend_n_367;
  wire frontend_n_368;
  wire frontend_n_369;
  wire frontend_n_370;
  wire frontend_n_371;
  wire frontend_n_372;
  wire frontend_n_373;
  wire frontend_n_374;
  wire frontend_n_375;
  wire frontend_n_376;
  wire frontend_n_378;
  wire frontend_n_386;
  wire frontend_n_387;
  wire frontend_n_388;
  wire frontend_n_389;
  wire frontend_n_390;
  wire frontend_n_391;
  wire frontend_n_392;
  wire frontend_n_393;
  wire frontend_n_395;
  wire frontend_n_396;
  wire frontend_n_402;
  wire frontend_n_403;
  wire frontend_n_404;
  wire frontend_n_409;
  wire frontend_n_410;
  wire frontend_n_416;
  wire frontend_n_419;
  wire frontend_n_44;
  wire frontend_n_49;
  wire frontend_n_51;
  wire frontend_n_52;
  wire frontend_n_54;
  wire frontend_n_92;
  wire got_e_reg;
  wire got_e_reg_0;
  wire host_clk;
  wire [4:4]\ibuf/_T_100 ;
  wire [15:0]\ibuf/_T_74 ;
  wire [1:1]\ibuf/_T_81 ;
  wire \ibuf/buf__pc ;
  wire \ibuf/buf__replay ;
  wire \ibuf/buf__xcpt_ae_inst ;
  wire [4:0]ibuf_io_inst_0_bits_inst_rd;
  wire [4:0]ibuf_io_inst_0_bits_inst_rs1;
  wire [4:0]ibuf_io_inst_0_bits_inst_rs2;
  wire [29:0]ibuf_io_inst_0_bits_raw;
  wire ibuf_io_inst_0_bits_xcpt0_ae_inst;
  wire [39:5]ibuf_io_pc;
  wire [0:0]\icache/_T_191_reg__0 ;
  wire \icache/invalidated ;
  wire \icache/load ;
  wire [0:0]\icache/p_0_in ;
  wire [8:0]\icache/p_0_in__0 ;
  wire \icache/p_12_in ;
  wire \icache/refill_one_beat ;
  wire \icache/refill_valid ;
  wire id_ctrl_alu_dw;
  wire [3:0]id_ctrl_alu_fn;
  wire id_ctrl_fence_i;
  wire id_ctrl_jal;
  wire id_ctrl_mem;
  wire [3:0]id_ctrl_mem_cmd;
  wire id_ctrl_rxs2;
  wire [1:0]id_ctrl_sel_alu1;
  wire [2:0]id_ctrl_sel_imm;
  wire id_ctrl_wxd;
  wire invalid_paddr;
  wire [25:0]io_enq_bits_address;
  wire [63:0]io_enq_bits_data;
  wire [1:0]io_enq_bits_param;
  wire [1:0]io_enq_bits_source;
  wire maybe_full_reg;
  wire maybe_full_reg_0;
  wire maybe_full_reg_1;
  wire mem_br_taken__reg_i_3_n_3;
  wire mem_br_taken__reg_i_4_n_0;
  wire mem_br_taken__reg_i_4_n_1;
  wire mem_br_taken__reg_i_4_n_2;
  wire mem_br_taken__reg_i_4_n_3;
  wire mem_br_taken__reg_i_6_n_0;
  wire mem_br_taken__reg_i_6_n_1;
  wire mem_br_taken__reg_i_6_n_2;
  wire mem_br_taken__reg_i_6_n_3;
  wire mem_br_taken__reg_i_7_n_0;
  wire mem_br_taken__reg_i_7_n_1;
  wire mem_br_taken__reg_i_7_n_2;
  wire mem_br_taken__reg_i_7_n_3;
  wire mem_br_taken__reg_i_8_n_0;
  wire mem_br_taken__reg_i_8_n_1;
  wire mem_br_taken__reg_i_8_n_2;
  wire mem_br_taken__reg_i_8_n_3;
  wire mem_br_taken__reg_i_9_n_0;
  wire mem_br_taken__reg_i_9_n_1;
  wire mem_br_taken__reg_i_9_n_2;
  wire mem_br_taken__reg_i_9_n_3;
  wire mem_ctrl_branch;
  wire mem_ctrl_fp;
  wire mem_ctrl_jal;
  wire mem_ctrl_jalr;
  wire mem_ctrl_mem;
  wire [3:2]mem_reg_cause;
  wire mem_reg_flush_pipe;
  wire [39:1]mem_reg_pc;
  wire mem_reg_replay_reg;
  wire [57:1]mem_reg_rs2;
  wire [57:41]mem_reg_rs20_in;
  wire mem_reg_rvc;
  wire mem_reg_sfence;
  wire mem_reg_slow_bypass;
  wire mem_reg_valid;
  wire mem_reg_xcpt;
  wire mem_reg_xcpt0;
  wire mem_reg_xcpt_interrupt;
  wire [4:0]mem_waddr;
  wire [39:0]p_0_in;
  wire [0:0]p_0_in_5;
  wire [29:0]p_1_in;
  wire p_31_in;
  wire p_4_in;
  wire pte_v;
  wire [19:0]ptw_io_dpath_ptbr_ppn;
  wire ptw_n_1;
  wire ptw_n_100;
  wire ptw_n_101;
  wire ptw_n_102;
  wire ptw_n_104;
  wire ptw_n_105;
  wire ptw_n_106;
  wire ptw_n_107;
  wire ptw_n_109;
  wire ptw_n_110;
  wire ptw_n_111;
  wire ptw_n_112;
  wire ptw_n_113;
  wire ptw_n_114;
  wire ptw_n_115;
  wire ptw_n_116;
  wire ptw_n_117;
  wire ptw_n_118;
  wire ptw_n_119;
  wire ptw_n_120;
  wire ptw_n_121;
  wire ptw_n_122;
  wire ptw_n_13;
  wire ptw_n_131;
  wire ptw_n_132;
  wire ptw_n_134;
  wire ptw_n_135;
  wire ptw_n_136;
  wire ptw_n_137;
  wire ptw_n_138;
  wire ptw_n_139;
  wire ptw_n_14;
  wire ptw_n_140;
  wire ptw_n_141;
  wire ptw_n_142;
  wire ptw_n_143;
  wire ptw_n_144;
  wire ptw_n_145;
  wire ptw_n_146;
  wire ptw_n_147;
  wire ptw_n_148;
  wire ptw_n_149;
  wire ptw_n_15;
  wire ptw_n_150;
  wire ptw_n_151;
  wire ptw_n_152;
  wire ptw_n_153;
  wire ptw_n_154;
  wire ptw_n_155;
  wire ptw_n_156;
  wire ptw_n_157;
  wire ptw_n_158;
  wire ptw_n_159;
  wire ptw_n_16;
  wire ptw_n_160;
  wire ptw_n_161;
  wire ptw_n_162;
  wire ptw_n_163;
  wire ptw_n_164;
  wire ptw_n_165;
  wire ptw_n_166;
  wire ptw_n_167;
  wire ptw_n_168;
  wire ptw_n_169;
  wire ptw_n_170;
  wire ptw_n_171;
  wire ptw_n_172;
  wire ptw_n_173;
  wire ptw_n_174;
  wire ptw_n_175;
  wire ptw_n_176;
  wire ptw_n_177;
  wire ptw_n_178;
  wire ptw_n_179;
  wire ptw_n_180;
  wire ptw_n_181;
  wire ptw_n_182;
  wire ptw_n_183;
  wire ptw_n_184;
  wire ptw_n_185;
  wire ptw_n_186;
  wire ptw_n_187;
  wire ptw_n_188;
  wire ptw_n_189;
  wire ptw_n_190;
  wire ptw_n_191;
  wire ptw_n_192;
  wire ptw_n_193;
  wire ptw_n_195;
  wire ptw_n_196;
  wire ptw_n_197;
  wire ptw_n_2;
  wire ptw_n_37;
  wire ptw_n_49;
  wire ptw_n_50;
  wire ptw_n_51;
  wire ptw_n_52;
  wire ptw_n_53;
  wire ptw_n_55;
  wire ptw_n_56;
  wire ptw_n_66;
  wire ptw_n_67;
  wire ptw_n_68;
  wire ptw_n_69;
  wire ptw_n_70;
  wire ptw_n_72;
  wire ptw_n_73;
  wire ptw_n_76;
  wire ptw_n_77;
  wire ptw_n_82;
  wire ptw_n_83;
  wire ptw_n_85;
  wire ptw_n_86;
  wire ptw_n_87;
  wire ptw_n_88;
  wire ptw_n_89;
  wire ptw_n_90;
  wire ptw_n_91;
  wire ptw_n_92;
  wire ptw_n_93;
  wire ptw_n_94;
  wire ptw_n_95;
  wire ptw_n_96;
  wire ptw_n_97;
  wire ptw_n_98;
  wire ptw_n_99;
  wire [0:0]q_reg;
  wire r_pte_d;
  wire [31:0]ram_address__T_63_data;
  wire [63:0]ram_data__T_63_data;
  wire [63:0]\ram_data_reg[63] ;
  wire \ram_id_reg[0] ;
  wire \ram_id_reg[3] ;
  wire \ram_id_reg[4] ;
  wire \ram_id_reg[5] ;
  wire [7:0]ram_mask__T_63_data;
  wire [0:0]\ram_opcode_reg[1] ;
  wire [1:0]ram_source__T_63_data;
  wire \ram_strb_reg[0] ;
  wire \ram_strb_reg[0]_0 ;
  wire \ram_strb_reg[1] ;
  wire \ram_strb_reg[2] ;
  wire \ram_strb_reg[2]_0 ;
  wire \ram_strb_reg[3] ;
  wire \ram_strb_reg[4] ;
  wire \ram_strb_reg[4]_0 ;
  wire \ram_strb_reg[5] ;
  wire \ram_strb_reg[6] ;
  wire \ram_strb_reg[6]_0 ;
  wire \ram_strb_reg[7] ;
  wire \ram_user_reg[6] ;
  wire release_ack_wait30_out;
  wire \remainder[103]_i_13_n_0 ;
  wire \remainder[103]_i_14_n_0 ;
  wire [2:0]\remainder_reg[103] ;
  wire [3:0]\remainder_reg[107] ;
  wire [3:0]\remainder_reg[107]_0 ;
  wire [3:0]\remainder_reg[111] ;
  wire [3:0]\remainder_reg[111]_0 ;
  wire [3:0]\remainder_reg[115] ;
  wire [0:0]\remainder_reg[115]_0 ;
  wire [2:0]\remainder_reg[115]_1 ;
  wire [3:0]\remainder_reg[64] ;
  wire [3:0]\remainder_reg[64]_0 ;
  wire [2:0]\remainder_reg[64]_1 ;
  wire resp_send_reg;
  wire s0_clk_en;
  wire [39:2]s1_pc;
  wire \s1_pc_reg[39]_i_12_n_0 ;
  wire \s1_pc_reg[39]_i_12_n_1 ;
  wire \s1_pc_reg[39]_i_12_n_2 ;
  wire \s1_pc_reg[39]_i_12_n_3 ;
  wire \s1_pc_reg[39]_i_14_n_0 ;
  wire \s1_pc_reg[39]_i_14_n_1 ;
  wire \s1_pc_reg[39]_i_14_n_2 ;
  wire \s1_pc_reg[39]_i_14_n_3 ;
  wire \s1_pc_reg[39]_i_16_n_0 ;
  wire \s1_pc_reg[39]_i_16_n_1 ;
  wire \s1_pc_reg[39]_i_16_n_2 ;
  wire \s1_pc_reg[39]_i_16_n_3 ;
  wire \s1_pc_reg[39]_i_21_n_0 ;
  wire \s1_pc_reg[39]_i_21_n_1 ;
  wire \s1_pc_reg[39]_i_21_n_2 ;
  wire \s1_pc_reg[39]_i_21_n_3 ;
  wire s1_release_data_valid;
  wire \s1_req_addr_reg[39]_i_13_n_0 ;
  wire \s1_req_addr_reg[39]_i_13_n_1 ;
  wire \s1_req_addr_reg[39]_i_13_n_2 ;
  wire \s1_req_addr_reg[39]_i_13_n_3 ;
  wire \s1_req_addr_reg[39]_i_4_n_0 ;
  wire \s1_req_addr_reg[39]_i_4_n_1 ;
  wire \s1_req_addr_reg[39]_i_4_n_2 ;
  wire \s1_req_addr_reg[39]_i_4_n_3 ;
  wire \s1_req_addr_reg[39]_i_6_n_0 ;
  wire \s1_req_addr_reg[39]_i_6_n_1 ;
  wire \s1_req_addr_reg[39]_i_6_n_2 ;
  wire \s1_req_addr_reg[39]_i_6_n_3 ;
  wire \s1_req_addr_reg[39]_i_8_n_0 ;
  wire \s1_req_addr_reg[39]_i_8_n_1 ;
  wire \s1_req_addr_reg[39]_i_8_n_2 ;
  wire \s1_req_addr_reg[39]_i_8_n_3 ;
  wire s1_valid;
  wire [38:1]s2_pc;
  wire s2_release_data_valid0;
  wire s2_replay;
  wire s2_uncached;
  wire s2_valid_reg;
  wire \saved_address_reg[1] ;
  wire \saved_address_reg[1]_0 ;
  wire \saved_address_reg[7] ;
  wire \saved_address_reg[7]_0 ;
  wire \saved_address_reg[7]_1 ;
  wire \saved_address_reg[7]_2 ;
  wire \saved_address_reg[7]_3 ;
  wire \saved_address_reg[7]_4 ;
  wire [1:0]sbus_auto_coupler_from_port_named_blkdevcontroller_passthru_in_0_a_bits_address;
  wire [3:0]sbus_auto_coupler_from_port_named_blkdevcontroller_passthru_in_1_a_bits_address;
  wire [2:0]sbus_auto_coupler_from_port_named_serialadapter_passthru_in_a_bits_address;
  wire [0:0]sbus_auto_coupler_from_port_named_serialadapter_passthru_in_a_bits_opcode;
  wire [2:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_opcode;
  wire [2:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_param;
  wire [3:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_size;
  wire sbus_auto_coupler_from_tile_named_tile_fixer_in_a_ready;
  wire sbus_auto_coupler_from_tile_named_tile_fixer_in_a_valid;
  wire sbus_auto_coupler_from_tile_named_tile_fixer_in_b_valid;
  wire sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_error;
  wire [2:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_opcode;
  wire [2:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_sink;
  wire [3:0]sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_size;
  wire sbus_auto_coupler_from_tile_named_tile_fixer_in_d_ready;
  wire [1:0]sbus_auto_coupler_to_mbus_nodelay_out_a_bits_opcode;
  wire [2:0]sbus_auto_coupler_to_mbus_nodelay_out_c_bits_size;
  wire sbus_auto_coupler_to_mbus_nodelay_out_d_ready;
  wire [3:0]\sendaddr_reg[11] ;
  wire \source_reg[0] ;
  wire [1:0]\source_reg[1] ;
  wire \source_reg[4] ;
  wire \state_reg[0] ;
  wire \state_reg[0]_0 ;
  wire \state_reg[0]_1 ;
  wire \state_reg[0]_2 ;
  wire \state_reg[0]_3 ;
  wire sync_xing_n_207;
  wire sync_xing_n_208;
  wire sync_xing_n_209;
  wire sync_xing_n_210;
  wire sync_xing_n_212;
  wire sync_xing_n_213;
  wire sync_xing_n_214;
  wire sync_xing_n_215;
  wire sync_xing_n_216;
  wire sync_xing_n_217;
  wire sync_xing_n_218;
  wire sync_xing_n_22;
  wire sync_xing_n_220;
  wire sync_xing_n_32;
  wire sync_xing_n_33;
  wire sync_xing_n_34;
  wire sync_xing_n_35;
  wire sync_xing_n_350;
  wire sync_xing_n_352;
  wire sync_xing_n_354;
  wire sync_xing_n_355;
  wire sync_xing_n_356;
  wire sync_xing_n_357;
  wire sync_xing_n_358;
  wire sync_xing_n_359;
  wire sync_xing_n_365;
  wire sync_xing_n_366;
  wire sync_xing_n_39;
  wire sync_xing_n_40;
  wire sync_xing_n_41;
  wire sync_xing_n_42;
  wire sync_xing_n_43;
  wire sync_xing_n_44;
  wire sync_xing_n_45;
  wire sync_xing_n_46;
  wire sync_xing_n_47;
  wire sync_xing_n_48;
  wire sync_xing_n_49;
  wire sync_xing_n_50;
  wire sync_xing_n_51;
  wire sync_xing_n_54;
  wire sync_xing_n_55;
  wire sync_xing_n_56;
  wire sync_xing_n_57;
  wire sync_xing_n_58;
  wire sync_xing_n_59;
  wire sys_reset_reg;
  wire [2:0]system_bus_xbar_auto_out_3_a_bits_param;
  wire tag_array_0_reg_i_10__0;
  wire tag_array_0_reg_i_11__0;
  wire tag_array_0_reg_i_12__0;
  wire tag_array_0_reg_i_13__0;
  wire tag_array_0_reg_i_13__0_0;
  wire tag_array_0_reg_i_8__0;
  wire tag_array_0_reg_i_9__0;
  wire target_reset;
  wire tile_auto_int_sync_xing_sinklzy_in_0_sync_0;
  wire tile_auto_int_sync_xing_sinklzy_in_0_sync_1;
  wire tile_auto_int_sync_xing_sinklzy_in_1_sync_0;
  wire tile_auto_int_sync_xing_sinklzy_in_2_sync_0;
  wire [0:0]tlMasterXbar_auto_in_0_a_bits_size;
  wire [31:0]tlMasterXbar_auto_in_0_b_bits_address;
  wire [1:0]tlMasterXbar_auto_in_0_b_bits_param;
  wire [3:0]tlMasterXbar_auto_in_0_b_bits_size;
  wire [63:0]tlMasterXbar_auto_in_0_d_bits_data;
  wire tlMasterXbar_auto_in_0_d_bits_error;
  wire [0:0]tlMasterXbar_auto_in_0_d_bits_opcode;
  wire [3:1]tlMasterXbar_auto_in_0_d_bits_size;
  wire [31:6]tlMasterXbar_auto_in_1_a_bits_address;
  wire [31:6]tlMasterXbar_auto_out_a_bits_address;
  wire [7:0]tlMasterXbar_auto_out_a_bits_mask;
  wire [2:2]tlMasterXbar_auto_out_a_bits_opcode;
  wire [2:1]tlMasterXbar_auto_out_a_bits_size;
  wire [1:1]tlMasterXbar_auto_out_b_bits_source;
  wire [31:0]tlMasterXbar_auto_out_c_bits_address;
  wire [63:0]tlMasterXbar_auto_out_c_bits_data;
  wire [1:0]tlMasterXbar_auto_out_c_bits_opcode;
  wire [1:0]tlMasterXbar_auto_out_c_bits_size;
  wire [0:0]tlMasterXbar_auto_out_c_bits_source;
  wire tlMasterXbar_n_10;
  wire tlMasterXbar_n_2;
  wire tlMasterXbar_n_4;
  wire tlMasterXbar_n_5;
  wire tlMasterXbar_n_6;
  wire tlMasterXbar_n_7;
  wire [3:3]\tlb/_GEN_29 ;
  wire \tlb/_GEN_36 ;
  wire \tlb/_T_1081 ;
  wire [1:1]\tlb/_T_1432 ;
  wire \tlb/_T_194 ;
  wire [30:12]\tlb/_T_200__0 ;
  wire \tlb/_T_210 ;
  wire [31:31]\tlb/_T_382 ;
  wire [31:31]\tlb/_T_382_3 ;
  wire [28:25]\tlb/_T_382__0 ;
  wire \tlb/_T_384 ;
  wire \tlb/_T_392 ;
  wire [16:16]\tlb/_T_480 ;
  wire \tlb/_T_482 ;
  wire [13:13]\tlb/_T_726 ;
  wire \tlb/_T_728 ;
  wire \tlb/_T_815 ;
  wire \tlb/_T_928 ;
  wire \tlb/_T_936 ;
  wire \tlb/_T_943 ;
  wire \tlb/_T_943_4 ;
  wire \tlb/_T_946 ;
  wire \tlb/_T_949 ;
  wire \tlb/_T_952 ;
  wire \tlb/bad_va ;
  wire \tlb/entries_1_u ;
  wire \tlb/entries_2_sr ;
  wire \tlb/entries_2_sx ;
  wire \tlb/entries_2_u ;
  wire \tlb/entries_3_g ;
  wire \tlb/entries_3_sr ;
  wire \tlb/entries_3_sx ;
  wire \tlb/entries_3_u ;
  wire \tlb/entries_4_sr ;
  wire \tlb/entries_4_sx ;
  wire \tlb/entries_4_u ;
  wire \tlb/hitsVec_4 ;
  wire [19:0]\tlb/p_0_in ;
  wire [19:13]\tlb/p_0_in_1 ;
  wire \tlb/p_13_in ;
  wire \tlb/p_2_in ;
  wire \tlb/pmp/_T_125 ;
  wire \tlb/pmp/_T_161 ;
  wire \tlb/pmp/_T_197 ;
  wire \tlb/pmp/_T_201 ;
  wire \tlb/pmp/_T_233 ;
  wire \tlb/pmp/_T_269 ;
  wire \tlb/pmp/_T_328 ;
  wire \tlb/pmp/_T_455 ;
  wire \tlb/pmp/_T_53 ;
  wire \tlb/pmp/_T_58 ;
  wire \tlb/pmp/_T_582 ;
  wire \tlb/pmp/_T_709 ;
  wire \tlb/pmp/_T_74 ;
  wire \tlb/pmp/_T_836 ;
  wire \tlb/pmp/_T_89 ;
  wire \tlb/pmp/_T_94 ;
  wire [1:0]\tlb/state ;
  wire [1:0]\tlb/state_2 ;
  wire tlb_io_req_bits_sfence_bits_rs2;
  wire traverse;
  wire trigA;
  wire trigB;
  wire \trig_pc[11]_i_2_n_0 ;
  wire \trig_pc[11]_i_3_n_0 ;
  wire \trig_pc[11]_i_4_n_0 ;
  wire \trig_pc[11]_i_5_n_0 ;
  wire \trig_pc[15]_i_2_n_0 ;
  wire \trig_pc[15]_i_3_n_0 ;
  wire \trig_pc[15]_i_4_n_0 ;
  wire \trig_pc[15]_i_5_n_0 ;
  wire \trig_pc[19]_i_2_n_0 ;
  wire \trig_pc[19]_i_3_n_0 ;
  wire \trig_pc[19]_i_4_n_0 ;
  wire \trig_pc[19]_i_5_n_0 ;
  wire \trig_pc[23]_i_2_n_0 ;
  wire \trig_pc[23]_i_3_n_0 ;
  wire \trig_pc[23]_i_4_n_0 ;
  wire \trig_pc[23]_i_5_n_0 ;
  wire \trig_pc[27]_i_2_n_0 ;
  wire \trig_pc[27]_i_3_n_0 ;
  wire \trig_pc[27]_i_4_n_0 ;
  wire \trig_pc[27]_i_5_n_0 ;
  wire \trig_pc[31]_i_2_n_0 ;
  wire \trig_pc[31]_i_3_n_0 ;
  wire \trig_pc[31]_i_4_n_0 ;
  wire \trig_pc[31]_i_5_n_0 ;
  wire \trig_pc[35]_i_2_n_0 ;
  wire \trig_pc[35]_i_3_n_0 ;
  wire \trig_pc[35]_i_4_n_0 ;
  wire \trig_pc[35]_i_5_n_0 ;
  wire \trig_pc[39]_i_2_n_0 ;
  wire \trig_pc[39]_i_3_n_0 ;
  wire \trig_pc[39]_i_4_n_0 ;
  wire \trig_pc[39]_i_5_n_0 ;
  wire \trig_pc[3]_i_2_n_0 ;
  wire \trig_pc[3]_i_3_n_0 ;
  wire \trig_pc[3]_i_4_n_0 ;
  wire \trig_pc[43]_i_2_n_0 ;
  wire \trig_pc[43]_i_3_n_0 ;
  wire \trig_pc[43]_i_4_n_0 ;
  wire \trig_pc[43]_i_5_n_0 ;
  wire \trig_pc[47]_i_2_n_0 ;
  wire \trig_pc[47]_i_3_n_0 ;
  wire \trig_pc[47]_i_4_n_0 ;
  wire \trig_pc[47]_i_5_n_0 ;
  wire \trig_pc[51]_i_2_n_0 ;
  wire \trig_pc[51]_i_3_n_0 ;
  wire \trig_pc[51]_i_4_n_0 ;
  wire \trig_pc[51]_i_5_n_0 ;
  wire \trig_pc[55]_i_2_n_0 ;
  wire \trig_pc[55]_i_3_n_0 ;
  wire \trig_pc[55]_i_4_n_0 ;
  wire \trig_pc[55]_i_5_n_0 ;
  wire \trig_pc[59]_i_2_n_0 ;
  wire \trig_pc[59]_i_3_n_0 ;
  wire \trig_pc[59]_i_4_n_0 ;
  wire \trig_pc[59]_i_5_n_0 ;
  wire \trig_pc[63]_i_4_n_0 ;
  wire \trig_pc[63]_i_5_n_0 ;
  wire \trig_pc[63]_i_6_n_0 ;
  wire \trig_pc[63]_i_7_n_0 ;
  wire \trig_pc[7]_i_2_n_0 ;
  wire \trig_pc[7]_i_3_n_0 ;
  wire \trig_pc[7]_i_4_n_0 ;
  wire \trig_pc[7]_i_5_n_0 ;
  wire \trig_pc_reg[11]_i_1_n_0 ;
  wire \trig_pc_reg[11]_i_1_n_1 ;
  wire \trig_pc_reg[11]_i_1_n_2 ;
  wire \trig_pc_reg[11]_i_1_n_3 ;
  wire \trig_pc_reg[11]_i_1_n_4 ;
  wire \trig_pc_reg[11]_i_1_n_5 ;
  wire \trig_pc_reg[11]_i_1_n_6 ;
  wire \trig_pc_reg[11]_i_1_n_7 ;
  wire \trig_pc_reg[15]_i_1_n_0 ;
  wire \trig_pc_reg[15]_i_1_n_1 ;
  wire \trig_pc_reg[15]_i_1_n_2 ;
  wire \trig_pc_reg[15]_i_1_n_3 ;
  wire \trig_pc_reg[15]_i_1_n_4 ;
  wire \trig_pc_reg[15]_i_1_n_5 ;
  wire \trig_pc_reg[15]_i_1_n_6 ;
  wire \trig_pc_reg[15]_i_1_n_7 ;
  wire \trig_pc_reg[19]_i_1_n_0 ;
  wire \trig_pc_reg[19]_i_1_n_1 ;
  wire \trig_pc_reg[19]_i_1_n_2 ;
  wire \trig_pc_reg[19]_i_1_n_3 ;
  wire \trig_pc_reg[19]_i_1_n_4 ;
  wire \trig_pc_reg[19]_i_1_n_5 ;
  wire \trig_pc_reg[19]_i_1_n_6 ;
  wire \trig_pc_reg[19]_i_1_n_7 ;
  wire \trig_pc_reg[23]_i_1_n_0 ;
  wire \trig_pc_reg[23]_i_1_n_1 ;
  wire \trig_pc_reg[23]_i_1_n_2 ;
  wire \trig_pc_reg[23]_i_1_n_3 ;
  wire \trig_pc_reg[23]_i_1_n_4 ;
  wire \trig_pc_reg[23]_i_1_n_5 ;
  wire \trig_pc_reg[23]_i_1_n_6 ;
  wire \trig_pc_reg[23]_i_1_n_7 ;
  wire \trig_pc_reg[27]_i_1_n_0 ;
  wire \trig_pc_reg[27]_i_1_n_1 ;
  wire \trig_pc_reg[27]_i_1_n_2 ;
  wire \trig_pc_reg[27]_i_1_n_3 ;
  wire \trig_pc_reg[27]_i_1_n_4 ;
  wire \trig_pc_reg[27]_i_1_n_5 ;
  wire \trig_pc_reg[27]_i_1_n_6 ;
  wire \trig_pc_reg[27]_i_1_n_7 ;
  wire \trig_pc_reg[31]_i_1_n_0 ;
  wire \trig_pc_reg[31]_i_1_n_1 ;
  wire \trig_pc_reg[31]_i_1_n_2 ;
  wire \trig_pc_reg[31]_i_1_n_3 ;
  wire \trig_pc_reg[31]_i_1_n_4 ;
  wire \trig_pc_reg[31]_i_1_n_5 ;
  wire \trig_pc_reg[31]_i_1_n_6 ;
  wire \trig_pc_reg[31]_i_1_n_7 ;
  wire \trig_pc_reg[35]_i_1_n_0 ;
  wire \trig_pc_reg[35]_i_1_n_1 ;
  wire \trig_pc_reg[35]_i_1_n_2 ;
  wire \trig_pc_reg[35]_i_1_n_3 ;
  wire \trig_pc_reg[35]_i_1_n_4 ;
  wire \trig_pc_reg[35]_i_1_n_5 ;
  wire \trig_pc_reg[35]_i_1_n_6 ;
  wire \trig_pc_reg[35]_i_1_n_7 ;
  wire \trig_pc_reg[39]_i_1_n_0 ;
  wire \trig_pc_reg[39]_i_1_n_1 ;
  wire \trig_pc_reg[39]_i_1_n_2 ;
  wire \trig_pc_reg[39]_i_1_n_3 ;
  wire \trig_pc_reg[39]_i_1_n_4 ;
  wire \trig_pc_reg[39]_i_1_n_5 ;
  wire \trig_pc_reg[39]_i_1_n_6 ;
  wire \trig_pc_reg[39]_i_1_n_7 ;
  wire \trig_pc_reg[3]_i_1_n_0 ;
  wire \trig_pc_reg[3]_i_1_n_1 ;
  wire \trig_pc_reg[3]_i_1_n_2 ;
  wire \trig_pc_reg[3]_i_1_n_3 ;
  wire \trig_pc_reg[3]_i_1_n_4 ;
  wire \trig_pc_reg[3]_i_1_n_5 ;
  wire \trig_pc_reg[3]_i_1_n_6 ;
  wire \trig_pc_reg[3]_i_1_n_7 ;
  wire \trig_pc_reg[43]_i_1_n_0 ;
  wire \trig_pc_reg[43]_i_1_n_1 ;
  wire \trig_pc_reg[43]_i_1_n_2 ;
  wire \trig_pc_reg[43]_i_1_n_3 ;
  wire \trig_pc_reg[43]_i_1_n_4 ;
  wire \trig_pc_reg[43]_i_1_n_5 ;
  wire \trig_pc_reg[43]_i_1_n_6 ;
  wire \trig_pc_reg[43]_i_1_n_7 ;
  wire \trig_pc_reg[47]_i_1_n_0 ;
  wire \trig_pc_reg[47]_i_1_n_1 ;
  wire \trig_pc_reg[47]_i_1_n_2 ;
  wire \trig_pc_reg[47]_i_1_n_3 ;
  wire \trig_pc_reg[47]_i_1_n_4 ;
  wire \trig_pc_reg[47]_i_1_n_5 ;
  wire \trig_pc_reg[47]_i_1_n_6 ;
  wire \trig_pc_reg[47]_i_1_n_7 ;
  wire \trig_pc_reg[51]_i_1_n_0 ;
  wire \trig_pc_reg[51]_i_1_n_1 ;
  wire \trig_pc_reg[51]_i_1_n_2 ;
  wire \trig_pc_reg[51]_i_1_n_3 ;
  wire \trig_pc_reg[51]_i_1_n_4 ;
  wire \trig_pc_reg[51]_i_1_n_5 ;
  wire \trig_pc_reg[51]_i_1_n_6 ;
  wire \trig_pc_reg[51]_i_1_n_7 ;
  wire \trig_pc_reg[55]_i_1_n_0 ;
  wire \trig_pc_reg[55]_i_1_n_1 ;
  wire \trig_pc_reg[55]_i_1_n_2 ;
  wire \trig_pc_reg[55]_i_1_n_3 ;
  wire \trig_pc_reg[55]_i_1_n_4 ;
  wire \trig_pc_reg[55]_i_1_n_5 ;
  wire \trig_pc_reg[55]_i_1_n_6 ;
  wire \trig_pc_reg[55]_i_1_n_7 ;
  wire \trig_pc_reg[59]_i_1_n_0 ;
  wire \trig_pc_reg[59]_i_1_n_1 ;
  wire \trig_pc_reg[59]_i_1_n_2 ;
  wire \trig_pc_reg[59]_i_1_n_3 ;
  wire \trig_pc_reg[59]_i_1_n_4 ;
  wire \trig_pc_reg[59]_i_1_n_5 ;
  wire \trig_pc_reg[59]_i_1_n_6 ;
  wire \trig_pc_reg[59]_i_1_n_7 ;
  wire \trig_pc_reg[63]_i_10_n_0 ;
  wire \trig_pc_reg[63]_i_10_n_1 ;
  wire \trig_pc_reg[63]_i_10_n_2 ;
  wire \trig_pc_reg[63]_i_10_n_3 ;
  wire \trig_pc_reg[63]_i_15_n_0 ;
  wire \trig_pc_reg[63]_i_15_n_1 ;
  wire \trig_pc_reg[63]_i_15_n_2 ;
  wire \trig_pc_reg[63]_i_15_n_3 ;
  wire \trig_pc_reg[63]_i_20_n_0 ;
  wire \trig_pc_reg[63]_i_20_n_1 ;
  wire \trig_pc_reg[63]_i_20_n_2 ;
  wire \trig_pc_reg[63]_i_20_n_3 ;
  wire \trig_pc_reg[63]_i_25_n_0 ;
  wire \trig_pc_reg[63]_i_25_n_1 ;
  wire \trig_pc_reg[63]_i_25_n_2 ;
  wire \trig_pc_reg[63]_i_25_n_3 ;
  wire \trig_pc_reg[63]_i_2_n_1 ;
  wire \trig_pc_reg[63]_i_2_n_2 ;
  wire \trig_pc_reg[63]_i_2_n_3 ;
  wire \trig_pc_reg[63]_i_2_n_4 ;
  wire \trig_pc_reg[63]_i_2_n_5 ;
  wire \trig_pc_reg[63]_i_2_n_6 ;
  wire \trig_pc_reg[63]_i_2_n_7 ;
  wire \trig_pc_reg[63]_i_3_n_3 ;
  wire \trig_pc_reg[63]_i_8_n_0 ;
  wire \trig_pc_reg[63]_i_8_n_1 ;
  wire \trig_pc_reg[63]_i_8_n_2 ;
  wire \trig_pc_reg[63]_i_8_n_3 ;
  wire \trig_pc_reg[7]_i_1_n_0 ;
  wire \trig_pc_reg[7]_i_1_n_1 ;
  wire \trig_pc_reg[7]_i_1_n_2 ;
  wire \trig_pc_reg[7]_i_1_n_3 ;
  wire \trig_pc_reg[7]_i_1_n_4 ;
  wire \trig_pc_reg[7]_i_1_n_5 ;
  wire \trig_pc_reg[7]_i_1_n_6 ;
  wire \trig_pc_reg[7]_i_1_n_7 ;
  wire \trig_state_reg[1]_i_12_n_0 ;
  wire \trig_state_reg[1]_i_12_n_1 ;
  wire \trig_state_reg[1]_i_12_n_2 ;
  wire \trig_state_reg[1]_i_12_n_3 ;
  wire \trig_state_reg[1]_i_17_n_0 ;
  wire \trig_state_reg[1]_i_17_n_1 ;
  wire \trig_state_reg[1]_i_17_n_2 ;
  wire \trig_state_reg[1]_i_17_n_3 ;
  wire \trig_state_reg[1]_i_22_n_0 ;
  wire \trig_state_reg[1]_i_22_n_1 ;
  wire \trig_state_reg[1]_i_22_n_2 ;
  wire \trig_state_reg[1]_i_22_n_3 ;
  wire \trig_state_reg[1]_i_3_n_3 ;
  wire \trig_state_reg[1]_i_5_n_0 ;
  wire \trig_state_reg[1]_i_5_n_1 ;
  wire \trig_state_reg[1]_i_5_n_2 ;
  wire \trig_state_reg[1]_i_5_n_3 ;
  wire \trig_state_reg[1]_i_7_n_0 ;
  wire \trig_state_reg[1]_i_7_n_1 ;
  wire \trig_state_reg[1]_i_7_n_2 ;
  wire \trig_state_reg[1]_i_7_n_3 ;
  wire value_1_reg;
  wire \value_1_reg[0] ;
  wire \value_1_reg[1] ;
  wire value_reg;
  wire value_reg_0;
  wire [2:0]wb_ctrl_csr;
  wire wb_ctrl_div;
  wire wb_ctrl_mem;
  wire wb_ctrl_wxd;
  wire [2:2]wb_reg_cause;
  wire [39:1]wb_reg_pc;
  wire wb_reg_replay;
  wire wb_reg_valid;
  wire wb_reg_xcpt;
  wire [4:0]wb_waddr;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h6)) 
    \bypass_mux_1[3]_i_7 
       (.I0(core_n_1782),
        .I1(ex_ctrl_alu_fn),
        .O(\bypass_mux_1[3]_i_7_n_0 ));
  CARRY4 \bypass_mux_1_reg[11]_i_2 
       (.CI(\bypass_mux_1_reg[7]_i_2_n_0 ),
        .CO({\bypass_mux_1_reg[11]_i_2_n_0 ,\bypass_mux_1_reg[11]_i_2_n_1 ,\bypass_mux_1_reg[11]_i_2_n_2 ,\bypass_mux_1_reg[11]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[11:8]),
        .O(dcacheArb_io_requestor_1_req_bits_addr[11:8]),
        .S({core_rep__5_n_0,core__271_n_0,core__270_n_0,core__269_n_0}));
  CARRY4 \bypass_mux_1_reg[15]_i_2 
       (.CI(\bypass_mux_1_reg[11]_i_2_n_0 ),
        .CO({\bypass_mux_1_reg[15]_i_2_n_0 ,\bypass_mux_1_reg[15]_i_2_n_1 ,\bypass_mux_1_reg[15]_i_2_n_2 ,\bypass_mux_1_reg[15]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[15:12]),
        .O(dcacheArb_io_requestor_1_req_bits_addr[15:12]),
        .S({core_rep__7_n_0,core__273_n_0,core__272_n_0,core_rep__6_n_0}));
  CARRY4 \bypass_mux_1_reg[19]_i_2 
       (.CI(\bypass_mux_1_reg[15]_i_2_n_0 ),
        .CO({\bypass_mux_1_reg[19]_i_2_n_0 ,\bypass_mux_1_reg[19]_i_2_n_1 ,\bypass_mux_1_reg[19]_i_2_n_2 ,\bypass_mux_1_reg[19]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[19:16]),
        .O(dcacheArb_io_requestor_1_req_bits_addr[19:16]),
        .S({core__276_n_0,core_rep__8_n_0,core__275_n_0,core__274_n_0}));
  CARRY4 \bypass_mux_1_reg[23]_i_2 
       (.CI(\bypass_mux_1_reg[19]_i_2_n_0 ),
        .CO({\bypass_mux_1_reg[23]_i_2_n_0 ,\bypass_mux_1_reg[23]_i_2_n_1 ,\bypass_mux_1_reg[23]_i_2_n_2 ,\bypass_mux_1_reg[23]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[23:20]),
        .O(dcacheArb_io_requestor_1_req_bits_addr[23:20]),
        .S({core__279_n_0,core__278_n_0,core_rep__9_n_0,core__277_n_0}));
  CARRY4 \bypass_mux_1_reg[27]_i_2 
       (.CI(\bypass_mux_1_reg[23]_i_2_n_0 ),
        .CO({\bypass_mux_1_reg[27]_i_2_n_0 ,\bypass_mux_1_reg[27]_i_2_n_1 ,\bypass_mux_1_reg[27]_i_2_n_2 ,\bypass_mux_1_reg[27]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[27:24]),
        .O(dcacheArb_io_requestor_1_req_bits_addr[27:24]),
        .S({core_rep__11_n_0,core__281_n_0,core__280_n_0,core_rep__10_n_0}));
  CARRY4 \bypass_mux_1_reg[3]_i_2 
       (.CI(\<const0> ),
        .CO({\bypass_mux_1_reg[3]_i_2_n_0 ,\bypass_mux_1_reg[3]_i_2_n_1 ,\bypass_mux_1_reg[3]_i_2_n_2 ,\bypass_mux_1_reg[3]_i_2_n_3 }),
        .CYINIT(core__320_n_0),
        .DI({alu_io_in1[3:1],core_n_1786}),
        .O(dcacheArb_io_requestor_1_req_bits_addr[3:0]),
        .S({core_rep__1_n_0,core_rep__0_n_0,core_rep_n_0,\bypass_mux_1[3]_i_7_n_0 }));
  CARRY4 \bypass_mux_1_reg[7]_i_2 
       (.CI(\bypass_mux_1_reg[3]_i_2_n_0 ),
        .CO({\bypass_mux_1_reg[7]_i_2_n_0 ,\bypass_mux_1_reg[7]_i_2_n_1 ,\bypass_mux_1_reg[7]_i_2_n_2 ,\bypass_mux_1_reg[7]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[7:4]),
        .O(dcacheArb_io_requestor_1_req_bits_addr[7:4]),
        .S({core__268_n_0,core_rep__4_n_0,core_rep__3_n_0,core_rep__2_n_0}));
  LUT5 #(
    .INIT(32'h556AAA6A)) 
    \bypass_mux_2[11]_i_3 
       (.I0(mem_reg_pc[11]),
        .I1(core_n_1114),
        .I2(mem_ctrl_jal),
        .I3(core_n_1355),
        .I4(mem_waddr[0]),
        .O(\bypass_mux_2[11]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[11]_i_4 
       (.I0(mem_reg_pc[10]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(core_n_1104),
        .O(\bypass_mux_2[11]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[11]_i_5 
       (.I0(mem_reg_pc[9]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(core_n_1105),
        .O(\bypass_mux_2[11]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[11]_i_6 
       (.I0(mem_reg_pc[8]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(core_n_1106),
        .O(\bypass_mux_2[11]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h556AAA6A)) 
    \bypass_mux_2[15]_i_3 
       (.I0(mem_reg_pc[15]),
        .I1(core_n_1119),
        .I2(mem_ctrl_jal),
        .I3(core_n_1355),
        .I4(_T_20810),
        .O(\bypass_mux_2[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h556AAA6A)) 
    \bypass_mux_2[15]_i_4 
       (.I0(mem_reg_pc[14]),
        .I1(core_n_1120),
        .I2(mem_ctrl_jal),
        .I3(core_n_1355),
        .I4(_T_20810),
        .O(\bypass_mux_2[15]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h556AAA6A)) 
    \bypass_mux_2[15]_i_5 
       (.I0(mem_reg_pc[13]),
        .I1(core_n_1121),
        .I2(mem_ctrl_jal),
        .I3(core_n_1355),
        .I4(_T_20810),
        .O(\bypass_mux_2[15]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h556AAA6A)) 
    \bypass_mux_2[15]_i_6 
       (.I0(mem_reg_pc[12]),
        .I1(core_n_1122),
        .I2(mem_ctrl_jal),
        .I3(core_n_1355),
        .I4(_T_20810),
        .O(\bypass_mux_2[15]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h556AAA6A)) 
    \bypass_mux_2[19]_i_3 
       (.I0(mem_reg_pc[19]),
        .I1(core_n_1115),
        .I2(mem_ctrl_jal),
        .I3(core_n_1355),
        .I4(_T_20810),
        .O(\bypass_mux_2[19]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h556AAA6A)) 
    \bypass_mux_2[19]_i_4 
       (.I0(mem_reg_pc[18]),
        .I1(core_n_1116),
        .I2(mem_ctrl_jal),
        .I3(core_n_1355),
        .I4(_T_20810),
        .O(\bypass_mux_2[19]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h556AAA6A)) 
    \bypass_mux_2[19]_i_5 
       (.I0(mem_reg_pc[17]),
        .I1(core_n_1117),
        .I2(mem_ctrl_jal),
        .I3(core_n_1355),
        .I4(_T_20810),
        .O(\bypass_mux_2[19]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h556AAA6A)) 
    \bypass_mux_2[19]_i_6 
       (.I0(mem_reg_pc[16]),
        .I1(core_n_1118),
        .I2(mem_ctrl_jal),
        .I3(core_n_1355),
        .I4(_T_20810),
        .O(\bypass_mux_2[19]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[23]_i_3 
       (.I0(mem_reg_pc[23]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(_T_20810),
        .O(\bypass_mux_2[23]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[23]_i_4 
       (.I0(mem_reg_pc[22]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(_T_20810),
        .O(\bypass_mux_2[23]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[23]_i_5 
       (.I0(mem_reg_pc[21]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(_T_20810),
        .O(\bypass_mux_2[23]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[23]_i_6 
       (.I0(mem_reg_pc[20]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(_T_20810),
        .O(\bypass_mux_2[23]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[27]_i_3 
       (.I0(mem_reg_pc[27]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(_T_20810),
        .O(\bypass_mux_2[27]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[27]_i_4 
       (.I0(mem_reg_pc[26]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(_T_20810),
        .O(\bypass_mux_2[27]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[27]_i_5 
       (.I0(mem_reg_pc[25]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(_T_20810),
        .O(\bypass_mux_2[27]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[27]_i_6 
       (.I0(mem_reg_pc[24]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(_T_20810),
        .O(\bypass_mux_2[27]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h1FE0)) 
    \bypass_mux_2[31]_i_4 
       (.I0(mem_ctrl_jal),
        .I1(core_n_1355),
        .I2(_T_20810),
        .I3(mem_reg_pc[31]),
        .O(\bypass_mux_2[31]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[31]_i_5 
       (.I0(mem_reg_pc[30]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(_T_20810),
        .O(\bypass_mux_2[31]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[31]_i_6 
       (.I0(mem_reg_pc[29]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(_T_20810),
        .O(\bypass_mux_2[31]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[31]_i_7 
       (.I0(mem_reg_pc[28]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(_T_20810),
        .O(\bypass_mux_2[31]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[7]_i_3 
       (.I0(mem_reg_pc[7]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(core_n_1107),
        .O(\bypass_mux_2[7]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[7]_i_4 
       (.I0(mem_reg_pc[6]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(core_n_1108),
        .O(\bypass_mux_2[7]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h56AA)) 
    \bypass_mux_2[7]_i_5 
       (.I0(mem_reg_pc[5]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1355),
        .I3(core_n_1109),
        .O(\bypass_mux_2[7]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h556AAA6A)) 
    \bypass_mux_2[7]_i_6 
       (.I0(mem_reg_pc[4]),
        .I1(core_n_1110),
        .I2(mem_ctrl_jal),
        .I3(core_n_1355),
        .I4(mem_waddr[4]),
        .O(\bypass_mux_2[7]_i_6_n_0 ));
  CARRY4 \bypass_mux_2_reg[11]_i_2 
       (.CI(\bypass_mux_2_reg[7]_i_2_n_0 ),
        .CO({\bypass_mux_2_reg[11]_i_2_n_0 ,\bypass_mux_2_reg[11]_i_2_n_1 ,\bypass_mux_2_reg[11]_i_2_n_2 ,\bypass_mux_2_reg[11]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(mem_reg_pc[11:8]),
        .O(p_0_in[11:8]),
        .S({\bypass_mux_2[11]_i_3_n_0 ,\bypass_mux_2[11]_i_4_n_0 ,\bypass_mux_2[11]_i_5_n_0 ,\bypass_mux_2[11]_i_6_n_0 }));
  CARRY4 \bypass_mux_2_reg[15]_i_2 
       (.CI(\bypass_mux_2_reg[11]_i_2_n_0 ),
        .CO({\bypass_mux_2_reg[15]_i_2_n_0 ,\bypass_mux_2_reg[15]_i_2_n_1 ,\bypass_mux_2_reg[15]_i_2_n_2 ,\bypass_mux_2_reg[15]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(mem_reg_pc[15:12]),
        .O(p_0_in[15:12]),
        .S({\bypass_mux_2[15]_i_3_n_0 ,\bypass_mux_2[15]_i_4_n_0 ,\bypass_mux_2[15]_i_5_n_0 ,\bypass_mux_2[15]_i_6_n_0 }));
  CARRY4 \bypass_mux_2_reg[19]_i_2 
       (.CI(\bypass_mux_2_reg[15]_i_2_n_0 ),
        .CO({\bypass_mux_2_reg[19]_i_2_n_0 ,\bypass_mux_2_reg[19]_i_2_n_1 ,\bypass_mux_2_reg[19]_i_2_n_2 ,\bypass_mux_2_reg[19]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(mem_reg_pc[19:16]),
        .O(p_0_in[19:16]),
        .S({\bypass_mux_2[19]_i_3_n_0 ,\bypass_mux_2[19]_i_4_n_0 ,\bypass_mux_2[19]_i_5_n_0 ,\bypass_mux_2[19]_i_6_n_0 }));
  CARRY4 \bypass_mux_2_reg[23]_i_2 
       (.CI(\bypass_mux_2_reg[19]_i_2_n_0 ),
        .CO({\bypass_mux_2_reg[23]_i_2_n_0 ,\bypass_mux_2_reg[23]_i_2_n_1 ,\bypass_mux_2_reg[23]_i_2_n_2 ,\bypass_mux_2_reg[23]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(mem_reg_pc[23:20]),
        .O(p_0_in[23:20]),
        .S({\bypass_mux_2[23]_i_3_n_0 ,\bypass_mux_2[23]_i_4_n_0 ,\bypass_mux_2[23]_i_5_n_0 ,\bypass_mux_2[23]_i_6_n_0 }));
  CARRY4 \bypass_mux_2_reg[27]_i_2 
       (.CI(\bypass_mux_2_reg[23]_i_2_n_0 ),
        .CO({\bypass_mux_2_reg[27]_i_2_n_0 ,\bypass_mux_2_reg[27]_i_2_n_1 ,\bypass_mux_2_reg[27]_i_2_n_2 ,\bypass_mux_2_reg[27]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(mem_reg_pc[27:24]),
        .O(p_0_in[27:24]),
        .S({\bypass_mux_2[27]_i_3_n_0 ,\bypass_mux_2[27]_i_4_n_0 ,\bypass_mux_2[27]_i_5_n_0 ,\bypass_mux_2[27]_i_6_n_0 }));
  CARRY4 \bypass_mux_2_reg[31]_i_2 
       (.CI(\bypass_mux_2_reg[27]_i_2_n_0 ),
        .CO({\bypass_mux_2_reg[31]_i_2_n_0 ,\bypass_mux_2_reg[31]_i_2_n_1 ,\bypass_mux_2_reg[31]_i_2_n_2 ,\bypass_mux_2_reg[31]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({_GEN_283,mem_reg_pc[30:28]}),
        .O(p_0_in[31:28]),
        .S({\bypass_mux_2[31]_i_4_n_0 ,\bypass_mux_2[31]_i_5_n_0 ,\bypass_mux_2[31]_i_6_n_0 ,\bypass_mux_2[31]_i_7_n_0 }));
  CARRY4 \bypass_mux_2_reg[35]_i_2 
       (.CI(\bypass_mux_2_reg[31]_i_2_n_0 ),
        .CO({\bypass_mux_2_reg[35]_i_2_n_0 ,\bypass_mux_2_reg[35]_i_2_n_1 ,\bypass_mux_2_reg[35]_i_2_n_2 ,\bypass_mux_2_reg[35]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({mem_reg_pc[34:32],core_n_1354}),
        .O(p_0_in[35:32]),
        .S({core__426_n_0,core__425_n_0,core__424_n_0,core__200_n_0}));
  CARRY4 \bypass_mux_2_reg[63]_i_3 
       (.CI(\bypass_mux_2_reg[35]_i_2_n_0 ),
        .CO({\bypass_mux_2_reg[63]_i_3_n_1 ,\bypass_mux_2_reg[63]_i_3_n_2 ,\bypass_mux_2_reg[63]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,mem_reg_pc[37:35]}),
        .O(p_0_in[39:36]),
        .S({core__429_n_0,core__430_n_0,core__428_n_0,core__427_n_0}));
  CARRY4 \bypass_mux_2_reg[7]_i_2 
       (.CI(core__201_i_1_n_0),
        .CO({\bypass_mux_2_reg[7]_i_2_n_0 ,\bypass_mux_2_reg[7]_i_2_n_1 ,\bypass_mux_2_reg[7]_i_2_n_2 ,\bypass_mux_2_reg[7]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(mem_reg_pc[7:4]),
        .O(p_0_in[7:4]),
        .S({\bypass_mux_2[7]_i_3_n_0 ,\bypass_mux_2[7]_i_4_n_0 ,\bypass_mux_2[7]_i_5_n_0 ,\bypass_mux_2[7]_i_6_n_0 }));
  Rocket core
       (.ADDRA(_T_1396__T_1415_addr),
        .CO(core_n_357),
        .D({core_n_91,core_n_92,core_n_93}),
        .DI({\remainder[103]_i_13_n_0 ,\remainder[103]_i_14_n_0 }),
        .E(core__185_n_0),
        .O(\div/_T_94 ),
        .Q(ex_ctrl_alu_fn),
        .S({core__420_n_0,core__421_n_0,core__422_n_0,core__423_n_0}),
        .SR(\icache/p_0_in ),
        ._GEN_274({_GEN_274[63:30],_GEN_274[9:0]}),
        ._T_100(\ibuf/_T_100 ),
        ._T_1005({_T_1005[6],_T_1005[4]}),
        ._T_1031(_T_1031[14]),
        ._T_1081(\tlb/_T_1081 ),
        ._T_1142({_T_1142[30],_T_1142[13:12]}),
        ._T_1156(_T_1156),
        ._T_121(\alu/_T_121 ),
        ._T_134(\bpu/_T_134 ),
        ._T_1406({_T_1406[63:2],_T_1406[0]}),
        ._T_1416(_T_1416),
        ._T_1432(\tlb/_T_1432 ),
        ._T_1573(_T_1573),
        ._T_1701(_T_1701[8:3]),
        ._T_1790(_T_1790),
        ._T_1821(_T_1821),
        ._T_1829(_T_1829),
        ._T_1844(_T_1844),
        .\_T_1883_reg[0] (core_n_1002),
        .\_T_1883_reg[1] (core_n_901),
        ._T_200__0({\tlb/_T_200__0 [30:29],\tlb/_T_200__0 [24:17],\tlb/_T_200__0 [15:14],\tlb/_T_200__0 [12]}),
        ._T_216(\div/_T_216 ),
        ._T_217(\alu/_T_217 ),
        .\_T_2547_reg[16]_0 (_T_2549),
        .\_T_2547_reg[16]_1 (frontend_n_403),
        .\_T_2547_reg[1]_0 (core_n_1095),
        .\_T_2547_reg[31]_0 (div_io_resp_bits_tag),
        .\_T_281_reg[0] (core__104_n_0),
        .\_T_281_reg[3] (\csr/_T_286__0 ),
        .\_T_294_reg[0] (core_n_894),
        .\_T_294_reg[0]_0 (core_n_997),
        .\_T_294_reg[0]_1 (core__103_n_0),
        .\_T_294_reg[3] (core_n_82),
        ._T_382(\tlb/_T_382 ),
        ._T_382_0(\tlb/_T_382_3 ),
        ._T_382__0({\tlb/_T_382__0 [28:27],\tlb/_T_382__0 [25]}),
        .\_T_389_reg[7] (core_n_1799),
        ._T_4068_ae_ld_reg(core_n_1837),
        ._T_4068_pf_ld_reg(core_n_1838),
        ._T_4068_pf_ld_reg_0(core_n_2079),
        ._T_4068_pf_ld_reg_1(core_n_2081),
        ._T_4068_pf_ld_reg_2(core_n_2082),
        ._T_4068_pf_ld_reg_3(core_n_2084),
        ._T_4068_pf_st_reg(core_n_2080),
        ._T_4068_pf_st_reg_0(core_n_2083),
        ._T_4068_pf_st_reg_1(core_n_2085),
        ._T_480(\tlb/_T_480 ),
        ._T_481(_T_481),
        ._T_4899(\csr/_T_4899 ),
        ._T_5044({\csr/_T_5044 [63],\csr/_T_5044 [4:0]}),
        ._T_5074(\csr/_T_5074 ),
        ._T_726(\tlb/_T_726 ),
        ._T_877(_T_877),
        ._T_889({_T_889[24:15],_T_889[11:7]}),
        ._T_909({_T_909[31],_T_909[29:26]}),
        ._T_931(_T_931),
        .\_T_973_reg[1] (core_n_1841),
        .\a_data_reg[63] (dcacheArb_io_requestor_1_s1_data_data),
        .alu_io_in1(alu_io_in1),
        .alu_io_in2({alu_io_in2[63:7],alu_io_in2[5:0]}),
        .bad_va(\tlb/bad_va ),
        .\buf__data_reg[12] (frontend_n_404),
        .\buf__data_reg[1] (core__55_n_0),
        .\buf__data_reg[1]_0 (core__51_n_0),
        .\buf__data_reg[1]_1 (core__699_n_0),
        .\buf__data_reg[1]_2 (core__704_n_0),
        .\buf__data_reg[1]_3 ({core__692_n_0,frontend_n_353}),
        .\buf__data_reg[2] (frontend_n_391),
        .\buf__data_reg[3] (frontend_n_358),
        .\buf__data_reg[3]_0 (core__695_n_0),
        .\buf__data_reg[3]_1 (id_ctrl_mem_cmd),
        .\buf__data_reg[3]_2 ({frontend_n_359,frontend_n_360}),
        .\buf__data_reg[3]_3 (id_ctrl_alu_fn),
        .\buf__data_reg[4] (frontend_n_372),
        .\buf__data_reg[4]_0 (frontend_n_392),
        .buf__pc(\ibuf/buf__pc ),
        .buf__replay(\ibuf/buf__replay ),
        .buf__xcpt_ae_inst(\ibuf/buf__xcpt_ae_inst ),
        .buf__xcpt_pf_inst_reg(frontend_n_355),
        .buf__xcpt_pf_inst_reg_0(core__95_n_0),
        .buf__xcpt_pf_inst_reg_1(frontend_n_354),
        .buf__xcpt_pf_inst_reg_2(core__96_n_0),
        .\bypass_mux_1_reg[0]_0 (core_n_1782),
        .\bypass_mux_1_reg[17]_0 (core_n_2302),
        .\bypass_mux_1_reg[18]_0 (core_n_2301),
        .\bypass_mux_1_reg[19]_0 (core_n_2300),
        .\bypass_mux_1_reg[1]_0 ({\alu/shin [63],\alu/shin [47],\alu/shin [31],\alu/shin [15]}),
        .\bypass_mux_1_reg[1]_1 (core_n_2315),
        .\bypass_mux_1_reg[1]_2 (core_n_2316),
        .\bypass_mux_1_reg[20]_0 (core_n_2299),
        .\bypass_mux_1_reg[21]_0 (core_n_2298),
        .\bypass_mux_1_reg[22]_0 (core_n_2297),
        .\bypass_mux_1_reg[23]_0 (core_n_2296),
        .\bypass_mux_1_reg[29]_0 (core_n_2285),
        .\bypass_mux_1_reg[29]_1 (core_n_2288),
        .\bypass_mux_1_reg[29]_2 (core_n_2293),
        .\bypass_mux_1_reg[29]_3 (core_n_2294),
        .\bypass_mux_1_reg[29]_4 (core_n_2295),
        .\bypass_mux_1_reg[2]_0 (core_n_2314),
        .\bypass_mux_1_reg[32]_0 (core_n_2203),
        .\bypass_mux_1_reg[33]_0 (core_n_2204),
        .\bypass_mux_1_reg[33]_1 (core_n_2284),
        .\bypass_mux_1_reg[33]_2 (core_n_2286),
        .\bypass_mux_1_reg[33]_3 (core_n_2291),
        .\bypass_mux_1_reg[33]_4 (core_n_2292),
        .\bypass_mux_1_reg[34]_0 (core_n_2205),
        .\bypass_mux_1_reg[34]_1 (core_n_2282),
        .\bypass_mux_1_reg[34]_2 (core_n_2283),
        .\bypass_mux_1_reg[34]_3 (core_n_2289),
        .\bypass_mux_1_reg[34]_4 (core_n_2290),
        .\bypass_mux_1_reg[35]_0 (core_n_2206),
        .\bypass_mux_1_reg[35]_1 (core_n_2280),
        .\bypass_mux_1_reg[35]_2 (core_n_2281),
        .\bypass_mux_1_reg[35]_3 (core_n_2287),
        .\bypass_mux_1_reg[36]_0 (core_n_2207),
        .\bypass_mux_1_reg[36]_1 (core_n_2279),
        .\bypass_mux_1_reg[36]_2 (\bpu/_T_66 ),
        .\bypass_mux_1_reg[37]_0 (core_n_2208),
        .\bypass_mux_1_reg[37]_1 (core_n_2277),
        .\bypass_mux_1_reg[37]_2 (core_n_2278),
        .\bypass_mux_1_reg[38]_0 (core_n_2209),
        .\bypass_mux_1_reg[38]_1 (core_n_2275),
        .\bypass_mux_1_reg[38]_2 (core_n_2276),
        .\bypass_mux_1_reg[38]_3 (\bpu/_T_39 ),
        .\bypass_mux_1_reg[39]_0 (core_n_2210),
        .\bypass_mux_1_reg[39]_1 (core_n_2273),
        .\bypass_mux_1_reg[39]_2 (core_n_2274),
        .\bypass_mux_1_reg[3]_0 (core_n_2313),
        .\bypass_mux_1_reg[40]_0 (core_n_2211),
        .\bypass_mux_1_reg[40]_1 (core_n_2271),
        .\bypass_mux_1_reg[40]_2 (core_n_2272),
        .\bypass_mux_1_reg[41]_0 (core_n_2212),
        .\bypass_mux_1_reg[41]_1 (core_n_2269),
        .\bypass_mux_1_reg[41]_2 (core_n_2270),
        .\bypass_mux_1_reg[42]_0 (core_n_2213),
        .\bypass_mux_1_reg[42]_1 (core_n_2267),
        .\bypass_mux_1_reg[42]_2 (core_n_2268),
        .\bypass_mux_1_reg[43]_0 (core_n_2214),
        .\bypass_mux_1_reg[43]_1 (core_n_2265),
        .\bypass_mux_1_reg[43]_2 (core_n_2266),
        .\bypass_mux_1_reg[44]_0 (core_n_2215),
        .\bypass_mux_1_reg[44]_1 (core_n_2263),
        .\bypass_mux_1_reg[44]_2 (core_n_2264),
        .\bypass_mux_1_reg[45]_0 (core_n_2216),
        .\bypass_mux_1_reg[45]_1 (core_n_2261),
        .\bypass_mux_1_reg[45]_2 (core_n_2262),
        .\bypass_mux_1_reg[46]_0 (core_n_2217),
        .\bypass_mux_1_reg[46]_1 (core_n_2259),
        .\bypass_mux_1_reg[46]_2 (core_n_2260),
        .\bypass_mux_1_reg[47]_0 (core_n_2218),
        .\bypass_mux_1_reg[47]_1 (core_n_2256),
        .\bypass_mux_1_reg[47]_2 (core_n_2257),
        .\bypass_mux_1_reg[48]_0 (core_n_2223),
        .\bypass_mux_1_reg[48]_1 (core_n_2254),
        .\bypass_mux_1_reg[48]_2 (core_n_2255),
        .\bypass_mux_1_reg[48]_3 (core_n_2318),
        .\bypass_mux_1_reg[49]_0 (core_n_2224),
        .\bypass_mux_1_reg[49]_1 (core_n_2253),
        .\bypass_mux_1_reg[49]_2 (core_n_2319),
        .\bypass_mux_1_reg[4]_0 (core_n_1777),
        .\bypass_mux_1_reg[50]_0 (core_n_2225),
        .\bypass_mux_1_reg[50]_1 (core_n_2252),
        .\bypass_mux_1_reg[50]_2 (core_n_2303),
        .\bypass_mux_1_reg[50]_3 (core_n_2320),
        .\bypass_mux_1_reg[51]_0 (core_n_2226),
        .\bypass_mux_1_reg[51]_1 (core_n_2251),
        .\bypass_mux_1_reg[51]_2 (core_n_2304),
        .\bypass_mux_1_reg[51]_3 (core_n_2321),
        .\bypass_mux_1_reg[52]_0 (core_n_2227),
        .\bypass_mux_1_reg[52]_1 (core_n_2250),
        .\bypass_mux_1_reg[52]_2 (core_n_2305),
        .\bypass_mux_1_reg[52]_3 (core_n_2322),
        .\bypass_mux_1_reg[53]_0 (core_n_2228),
        .\bypass_mux_1_reg[53]_1 (core_n_2249),
        .\bypass_mux_1_reg[53]_2 (core_n_2306),
        .\bypass_mux_1_reg[53]_3 (core_n_2323),
        .\bypass_mux_1_reg[54]_0 (core_n_2229),
        .\bypass_mux_1_reg[54]_1 (core_n_2248),
        .\bypass_mux_1_reg[54]_2 (core_n_2307),
        .\bypass_mux_1_reg[54]_3 (core_n_2324),
        .\bypass_mux_1_reg[55]_0 (core_n_2230),
        .\bypass_mux_1_reg[55]_1 (core_n_2247),
        .\bypass_mux_1_reg[55]_2 (core_n_2308),
        .\bypass_mux_1_reg[55]_3 (core_n_2325),
        .\bypass_mux_1_reg[56]_0 (core_n_2231),
        .\bypass_mux_1_reg[56]_1 (core_n_2246),
        .\bypass_mux_1_reg[56]_2 (core_n_2309),
        .\bypass_mux_1_reg[56]_3 (core_n_2326),
        .\bypass_mux_1_reg[57]_0 (core_n_2232),
        .\bypass_mux_1_reg[57]_1 (core_n_2245),
        .\bypass_mux_1_reg[57]_2 (core_n_2310),
        .\bypass_mux_1_reg[57]_3 (core_n_2327),
        .\bypass_mux_1_reg[58]_0 (core_n_2233),
        .\bypass_mux_1_reg[58]_1 (core_n_2244),
        .\bypass_mux_1_reg[58]_2 (core_n_2311),
        .\bypass_mux_1_reg[58]_3 (core_n_2328),
        .\bypass_mux_1_reg[59]_0 (core_n_2234),
        .\bypass_mux_1_reg[59]_1 (core_n_2243),
        .\bypass_mux_1_reg[59]_2 (core_n_2312),
        .\bypass_mux_1_reg[59]_3 (core_n_2329),
        .\bypass_mux_1_reg[60]_0 (core_n_2219),
        .\bypass_mux_1_reg[60]_1 (core_n_2242),
        .\bypass_mux_1_reg[61]_0 (core_n_2220),
        .\bypass_mux_1_reg[61]_1 (core_n_2241),
        .\bypass_mux_1_reg[62]_0 (core_n_2221),
        .\bypass_mux_1_reg[62]_1 (core_n_2240),
        .\bypass_mux_1_reg[63]_0 (core_n_2222),
        .\bypass_mux_1_reg[63]_1 (_T_2181),
        .\bypass_mux_1_reg[63]_2 (_T_2179),
        .\bypass_mux_1_reg[6]_0 (core_n_1776),
        .\bypass_mux_1_reg[6]_1 (ex_ctrl_sel_imm),
        .\bypass_mux_2_reg[31]_0 ({_GEN_283,mem_reg_pc[30:28]}),
        .\bypass_mux_2_reg[35]_0 (core_n_1355),
        .\bypass_mux_2_reg[38]_0 (core_n_1329),
        .\bypass_mux_2_reg[63]_0 (_T_2520),
        .\bypass_mux_2_reg[63]_1 (_T_2522),
        .\bypass_mux_2_reg[63]_2 ({core__7_n_0,core__8_n_0,core__9_n_0,core__10_n_0,core__11_n_0,core__12_n_0,core__13_n_0,core__14_n_0,core__15_n_0,core__16_n_0,core__17_n_0,core__18_n_0,core__19_n_0,core__20_n_0,core__21_n_0,core__22_n_0,core__23_n_0,core__24_n_0,core__25_n_0,core__26_n_0,core__27_n_0,core__28_n_0,core__29_n_0,core__30_n_0,core__31_n_0,core__32_n_0,core__33_n_0,core__34_n_0,core__35_n_0,core__36_n_0,core__37_n_0,core__38_n_0,p_1_in}),
        .\bypass_mux_2_reg[9]_0 (\div/p_1_in ),
        .\count_reg[0] (core_n_103),
        .\count_reg[1] (ptw_n_85),
        .\count_reg[1]_0 (ptw_n_90),
        .\count_reg[1]_1 (ptw_n_113),
        .\count_reg[1]_2 (ptw_n_118),
        .csr_io_bp_0_control_action(csr_io_bp_0_control_action),
        .csr_io_bp_0_control_m(csr_io_bp_0_control_m),
        .csr_io_bp_0_control_s(csr_io_bp_0_control_s),
        .csr_io_bp_0_control_u(csr_io_bp_0_control_u),
        .csr_io_status_debug(csr_io_status_debug),
        .csr_io_tval(csr_io_tval),
        .dcacheArb_io_requestor_1_ordered(dcacheArb_io_requestor_1_ordered),
        .dcacheArb_io_requestor_1_replay_next(dcacheArb_io_requestor_1_replay_next),
        .dcacheArb_io_requestor_1_req_bits_addr(dcacheArb_io_requestor_1_req_bits_addr[32:0]),
        .dcacheArb_io_requestor_1_req_bits_typ(dcacheArb_io_requestor_1_req_bits_typ),
        .dcacheArb_io_requestor_1_req_ready(dcacheArb_io_requestor_1_req_ready),
        .dcacheArb_io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),
        .dcacheArb_io_requestor_1_resp_bits_data({dcacheArb_io_requestor_1_resp_bits_data[63:30],dcacheArb_io_requestor_1_resp_bits_data[9:0]}),
        .dcacheArb_io_requestor_1_resp_bits_data_word_bypass(dcacheArb_io_requestor_1_resp_bits_data_word_bypass),
        .dcacheArb_io_requestor_1_resp_bits_replay(dcacheArb_io_requestor_1_resp_bits_replay),
        .dcacheArb_io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),
        .dcacheArb_io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),
        .dcacheArb_io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),
        .dcacheArb_io_requestor_1_s2_xcpt_ma_ld(dcacheArb_io_requestor_1_s2_xcpt_ma_ld),
        .dcacheArb_io_requestor_1_s2_xcpt_ma_st(dcacheArb_io_requestor_1_s2_xcpt_ma_st),
        .dcacheArb_io_requestor_1_s2_xcpt_pf_ld(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
        .dcacheArb_io_requestor_1_s2_xcpt_pf_st(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
        .dcache_io_cpu_invalidate_lr(dcache_io_cpu_invalidate_lr),
        .dcache_io_ptw_resp_bits_ae(dcache_io_ptw_resp_bits_ae),
        .dcache_io_ptw_resp_bits_homogeneous(dcache_io_ptw_resp_bits_homogeneous),
        .dcache_io_ptw_resp_bits_level(dcache_io_ptw_resp_bits_level),
        .dcache_io_ptw_resp_valid(dcache_io_ptw_resp_valid),
        .dcache_io_ptw_status_mxr(dcache_io_ptw_status_mxr),
        .dcache_io_ptw_status_sum(dcache_io_ptw_status_sum),
        .\divisor_reg[15] ({core__337_n_0,core__338_n_0,core__339_n_0}),
        .\divisor_reg[15]_0 ({core__333_n_0,core__334_n_0,core__335_n_0,core__336_n_0}),
        .\divisor_reg[15]_1 ({core__329_n_0,core__330_n_0,core__331_n_0,core__332_n_0}),
        .\divisor_reg[15]_2 ({core__325_n_0,core__326_n_0,core__327_n_0,core__328_n_0}),
        .\divisor_reg[15]_3 ({core_rep__24_n_0,core_rep__23_n_0,core__340_n_0,core__341_n_0}),
        .\divisor_reg[15]_4 ({core__342_i_20_n_0,core__342_i_21_n_0,core__342_i_22_n_0,core__342_i_23_n_0}),
        .\divisor_reg[15]_5 ({core_rep__28_n_0,core_rep__27_n_0,core_rep__26_n_0,core_rep__25_n_0}),
        .\divisor_reg[15]_6 ({core__342_i_12_n_0,core__342_i_13_n_0,core__342_i_14_n_0,core__342_i_15_n_0}),
        .\divisor_reg[15]_7 ({core_rep__32_n_0,core_rep__31_n_0,core_rep__30_n_0,core_rep__29_n_0}),
        .\divisor_reg[15]_8 ({core__342_i_4_n_0,core__342_i_5_n_0}),
        .\divisor_reg[18] (core__190_n_0),
        .\divisor_reg[1] (core__189_n_0),
        .\divisor_reg[32] ({core__342_i_6_n_0,core__459_n_0,core_rep__33_n_0}),
        .\divisor_reg[32]_0 ({core__349_n_0,core__350_n_0,core__351_n_0,core__352_n_0}),
        .\divisor_reg[32]_1 ({core__345_n_0,core__346_n_0,core__347_n_0,core__348_n_0}),
        .\divisor_reg[35] (core__187_n_0),
        .\divisor_reg[51] ({core__353_n_0,core__354_n_0,core__355_n_0,core__356_n_0}),
        .\divisor_reg[52] (core__188_n_0),
        .\divisor_reg[57] ({mem_reg_rs2[57],mem_reg_rs2[41],mem_reg_rs2[25],mem_reg_rs2[7:6],mem_reg_rs2[1]}),
        .doUncachedResp_reg(dcache_n_553),
        .\elts_0_data_reg[15] (\ibuf/_T_74 ),
        .\elts_0_pc_reg[38] (\bpu/_T_105 ),
        .\elts_0_pc_reg[39] ({ibuf_io_pc[39:37],ibuf_io_pc[35],ibuf_io_pc[33],ibuf_io_pc[31],ibuf_io_pc[29],ibuf_io_pc[27],ibuf_io_pc[25],ibuf_io_pc[23],ibuf_io_pc[21],ibuf_io_pc[19],ibuf_io_pc[17],ibuf_io_pc[15],ibuf_io_pc[13],ibuf_io_pc[11],ibuf_io_pc[9],ibuf_io_pc[7],ibuf_io_pc[5]}),
        .elts_0_xcpt_ae_inst_reg(frontend_n_419),
        .\ex_cause_reg[1]_0 (csr_io_bp_0_control_tmatch),
        .\ex_cause_reg[1]_1 (core_n_2102),
        .\ex_cause_reg[1]_10 ({core_n_2133,core_n_2134,core_n_2135,core_n_2136}),
        .\ex_cause_reg[1]_11 ({core_n_2137,core_n_2138,core_n_2139,core_n_2140}),
        .\ex_cause_reg[1]_12 ({core_n_2141,core_n_2142,core_n_2143,core_n_2144}),
        .\ex_cause_reg[1]_13 ({core_n_2145,core_n_2146,core_n_2147}),
        .\ex_cause_reg[1]_14 ({core_n_2148,core_n_2149,core_n_2150}),
        .\ex_cause_reg[1]_2 ({core_n_2103,core_n_2104,core_n_2105}),
        .\ex_cause_reg[1]_3 ({core_n_2106,core_n_2107,core_n_2108}),
        .\ex_cause_reg[1]_4 ({core_n_2109,core_n_2110,core_n_2111,core_n_2112}),
        .\ex_cause_reg[1]_5 ({core_n_2113,core_n_2114,core_n_2115,core_n_2116}),
        .\ex_cause_reg[1]_6 ({core_n_2117,core_n_2118,core_n_2119,core_n_2120}),
        .\ex_cause_reg[1]_7 ({core_n_2121,core_n_2122,core_n_2123,core_n_2124}),
        .\ex_cause_reg[1]_8 ({core_n_2125,core_n_2126,core_n_2127,core_n_2128}),
        .\ex_cause_reg[1]_9 ({core_n_2129,core_n_2130,core_n_2131,core_n_2132}),
        .ex_ctrl_alu_dw_reg_0(core__6_n_0),
        .ex_ctrl_alu_dw_reg_1(core__161_n_0),
        .ex_ctrl_alu_dw_reg_10(core__152_n_0),
        .ex_ctrl_alu_dw_reg_11(core__151_n_0),
        .ex_ctrl_alu_dw_reg_12(core__150_n_0),
        .ex_ctrl_alu_dw_reg_13(core__149_n_0),
        .ex_ctrl_alu_dw_reg_14(core__148_n_0),
        .ex_ctrl_alu_dw_reg_15(core__147_n_0),
        .ex_ctrl_alu_dw_reg_16(core__146_n_0),
        .ex_ctrl_alu_dw_reg_17(core__145_n_0),
        .ex_ctrl_alu_dw_reg_18(core__144_n_0),
        .ex_ctrl_alu_dw_reg_19(core__143_n_0),
        .ex_ctrl_alu_dw_reg_2(core__160_n_0),
        .ex_ctrl_alu_dw_reg_20(core__142_n_0),
        .ex_ctrl_alu_dw_reg_21(core__141_n_0),
        .ex_ctrl_alu_dw_reg_22(core__140_n_0),
        .ex_ctrl_alu_dw_reg_23(core__139_n_0),
        .ex_ctrl_alu_dw_reg_24(core__138_n_0),
        .ex_ctrl_alu_dw_reg_25(core__137_n_0),
        .ex_ctrl_alu_dw_reg_26(core__136_n_0),
        .ex_ctrl_alu_dw_reg_27(core__135_n_0),
        .ex_ctrl_alu_dw_reg_28(core__134_n_0),
        .ex_ctrl_alu_dw_reg_29(core__133_n_0),
        .ex_ctrl_alu_dw_reg_3(core__159_n_0),
        .ex_ctrl_alu_dw_reg_30(core__132_n_0),
        .ex_ctrl_alu_dw_reg_31(core__131_n_0),
        .ex_ctrl_alu_dw_reg_32(core__130_n_0),
        .ex_ctrl_alu_dw_reg_33(core__640_n_0),
        .ex_ctrl_alu_dw_reg_4(core__158_n_0),
        .ex_ctrl_alu_dw_reg_5(core__157_n_0),
        .ex_ctrl_alu_dw_reg_6(core__156_n_0),
        .ex_ctrl_alu_dw_reg_7(core__155_n_0),
        .ex_ctrl_alu_dw_reg_8(core__154_n_0),
        .ex_ctrl_alu_dw_reg_9(core__153_n_0),
        .\ex_ctrl_alu_fn_reg[3]_0 (core__441_n_0),
        .\ex_ctrl_alu_fn_reg[3]_1 (core__435_n_0),
        .\ex_ctrl_alu_fn_reg[3]_2 (core__437_n_0),
        .\ex_ctrl_alu_fn_reg[3]_3 (core__438_n_0),
        .\ex_ctrl_alu_fn_reg[3]_4 (core__439_n_0),
        .\ex_ctrl_alu_fn_reg[3]_5 (core__648_n_0),
        .\ex_ctrl_alu_fn_reg[3]_6 (core__662_n_0),
        .\ex_ctrl_alu_fn_reg[3]_7 (core__663_n_0),
        .\ex_ctrl_alu_fn_reg[3]_8 (core__284_n_0),
        .\ex_ctrl_alu_fn_reg[3]_9 (\alu/_T_31 ),
        .\ex_ctrl_csr_reg[0]_0 (frontend_n_225),
        .\ex_ctrl_csr_reg[1]_0 (frontend_n_231),
        .\ex_ctrl_csr_reg[2]_0 (core__715_n_0),
        .ex_ctrl_div(ex_ctrl_div),
        .ex_ctrl_div_reg_0(core__183_n_0),
        .ex_ctrl_fence_i(ex_ctrl_fence_i),
        .ex_ctrl_jalr(ex_ctrl_jalr),
        .ex_ctrl_mem_reg_0(core_n_1090),
        .ex_ctrl_mem_reg_1(core_n_1092),
        .ex_ctrl_mem_reg_10(core_n_1360),
        .ex_ctrl_mem_reg_11(core_n_1362),
        .ex_ctrl_mem_reg_2(core_n_1096),
        .ex_ctrl_mem_reg_3(core_n_1098),
        .ex_ctrl_mem_reg_4(core_n_1099),
        .ex_ctrl_mem_reg_5(core_n_1100),
        .ex_ctrl_mem_reg_6(core_n_1128),
        .ex_ctrl_mem_reg_7(core_n_1238),
        .ex_ctrl_mem_reg_8(core_n_1239),
        .ex_ctrl_mem_reg_9(core_n_1240),
        .\ex_ctrl_mem_type_reg[0]_0 ({mem_reg_rs20_in[57],mem_reg_rs20_in[41]}),
        .\ex_ctrl_sel_alu1_reg[0]_0 (core_n_1681),
        .\ex_ctrl_sel_alu1_reg[1]_0 (core_n_1680),
        .ex_ctrl_sel_alu2(ex_ctrl_sel_alu2),
        .\ex_ctrl_sel_alu2_reg[1]_0 (core_n_95),
        .\ex_ctrl_sel_alu2_reg[1]_1 (core_n_890),
        .\ex_ctrl_sel_alu2_reg[1]_2 (core_n_891),
        .\ex_ctrl_sel_alu2_reg[1]_3 (core_n_892),
        .\ex_ctrl_sel_alu2_reg[1]_4 (core_n_1089),
        .\ex_ctrl_sel_alu2_reg[1]_5 (core_n_1097),
        .\ex_ctrl_sel_imm_reg[1]_0 (core__321_n_0),
        .\ex_ctrl_sel_imm_reg[1]_1 (core__322_n_0),
        .ex_ctrl_wxd(ex_ctrl_wxd),
        .ex_ctrl_wxd_reg_0(core__706_n_0),
        .ex_ctrl_wxd_reg_1(ex_reg_rs_lsb_1),
        .ex_reg_flush_pipe(ex_reg_flush_pipe),
        .\ex_reg_inst_reg[10]_0 (frontend_n_373),
        .\ex_reg_inst_reg[10]_1 (core__639_n_0),
        .\ex_reg_inst_reg[10]_2 (core__641_n_0),
        .\ex_reg_inst_reg[10]_3 (core__643_n_0),
        .\ex_reg_inst_reg[10]_4 (core__644_n_0),
        .\ex_reg_inst_reg[10]_5 (core__646_n_0),
        .\ex_reg_inst_reg[10]_6 (core__645_n_0),
        .\ex_reg_inst_reg[10]_7 (core__647_n_0),
        .\ex_reg_inst_reg[11]_0 ({core_n_2086,core_n_2087,core_n_2088,core_n_2089,core_n_2090,core_n_2091,core_n_2092,core_n_2093,core_n_2094,core_n_2095,core_n_2096,core_n_2097,core_n_2098,core_n_2099,core_n_2100,core_n_2101}),
        .\ex_reg_inst_reg[26]_0 (core__440_n_0),
        .\ex_reg_pc_reg[39]_0 ({core_n_1069,core_n_1070,core_n_1071,core_n_1072,core_n_1073,core_n_1074,core_n_1075,core_n_1076,core_n_1077,core_n_1078,core_n_1079,core_n_1080,core_n_1081,core_n_1082,core_n_1083,core_n_1084,core_n_1085,core_n_1086,core_n_1087,core_n_1088}),
        .\ex_reg_pc_reg[39]_1 (core__157_i_3_n_4),
        .ex_reg_rs_bypass_0_reg_0(core_n_32),
        .ex_reg_rs_bypass_0_reg_1(core__4_n_0),
        .ex_reg_rs_bypass_1_reg_0(core_n_1093),
        .\ex_reg_rs_lsb_0_reg[0]_0 (core_n_1094),
        .\ex_reg_rs_lsb_0_reg[0]_1 (core_n_1102),
        .\ex_reg_rs_lsb_0_reg[1]_0 (core_n_1129),
        .\ex_reg_rs_msb_0_reg[10]_0 (core_n_1258),
        .\ex_reg_rs_msb_0_reg[11]_0 (core_n_1261),
        .\ex_reg_rs_msb_0_reg[12]_0 (core_n_1262),
        .\ex_reg_rs_msb_0_reg[13]_0 (core_n_1263),
        .\ex_reg_rs_msb_0_reg[14]_0 (core_n_1264),
        .\ex_reg_rs_msb_0_reg[15]_0 (core_n_1265),
        .\ex_reg_rs_msb_0_reg[16]_0 (core_n_1266),
        .\ex_reg_rs_msb_0_reg[17]_0 (core_n_1267),
        .\ex_reg_rs_msb_0_reg[18]_0 (core_n_1268),
        .\ex_reg_rs_msb_0_reg[19]_0 (core_n_1269),
        .\ex_reg_rs_msb_0_reg[20]_0 (core_n_1270),
        .\ex_reg_rs_msb_0_reg[21]_0 (core_n_1271),
        .\ex_reg_rs_msb_0_reg[22]_0 (core_n_1272),
        .\ex_reg_rs_msb_0_reg[23]_0 (core_n_1273),
        .\ex_reg_rs_msb_0_reg[24]_0 (core_n_1274),
        .\ex_reg_rs_msb_0_reg[25]_0 (core_n_1275),
        .\ex_reg_rs_msb_0_reg[26]_0 (core_n_1276),
        .\ex_reg_rs_msb_0_reg[27]_0 (div_io_resp_bits_data),
        .\ex_reg_rs_msb_0_reg[27]_1 (core_n_1277),
        .\ex_reg_rs_msb_0_reg[8]_0 (core_n_1259),
        .\ex_reg_rs_msb_0_reg[9]_0 (core_n_1260),
        .\ex_reg_rs_msb_1_reg[29]_0 ({\div/_GEN_36 ,\div/_GEN_35 [1],\div/_T_122 ,\div/_GEN_35 [0]}),
        .\ex_reg_rs_msb_1_reg[61]_0 (core_n_1249),
        .\ex_reg_rs_msb_1_reg[61]_1 (_T_1396__T_2475_addr),
        .\ex_reg_rs_msb_1_reg[61]_2 (core_n_1323),
        .ex_reg_rvc_reg_0(core_n_1256),
        .ex_reg_rvc_reg_1(core__5_n_0),
        .ex_reg_rvc_reg_10(core__655_n_0),
        .ex_reg_rvc_reg_11(core__656_n_0),
        .ex_reg_rvc_reg_12(core__657_n_0),
        .ex_reg_rvc_reg_13(core__658_n_0),
        .ex_reg_rvc_reg_14(core__659_n_0),
        .ex_reg_rvc_reg_15(core__660_n_0),
        .ex_reg_rvc_reg_16(core__661_n_0),
        .ex_reg_rvc_reg_2(core__638_n_0),
        .ex_reg_rvc_reg_3(core__642_n_0),
        .ex_reg_rvc_reg_4(core__649_n_0),
        .ex_reg_rvc_reg_5(core__650_n_0),
        .ex_reg_rvc_reg_6(core__651_n_0),
        .ex_reg_rvc_reg_7(core__652_n_0),
        .ex_reg_rvc_reg_8(core__653_n_0),
        .ex_reg_rvc_reg_9(core__654_n_0),
        .ex_reg_valid(ex_reg_valid),
        .ex_reg_xcpt(ex_reg_xcpt),
        .ex_reg_xcpt_interrupt(ex_reg_xcpt_interrupt),
        .ex_sfence(ex_sfence),
        .frontend_io_cpu_req_bits_speculative(frontend_io_cpu_req_bits_speculative),
        .frontend_io_cpu_resp_bits_data({frontend_io_cpu_resp_bits_data[28],frontend_io_cpu_resp_bits_data[12]}),
        .frontend_io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
        .frontend_io_cpu_resp_bits_replay(frontend_io_cpu_resp_bits_replay),
        .frontend_io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),
        .frontend_io_cpu_resp_bits_xcpt_pf_inst(frontend_io_cpu_resp_bits_xcpt_pf_inst),
        .frontend_io_cpu_resp_valid(frontend_io_cpu_resp_valid),
        .frontend_io_cpu_sfence_valid(frontend_io_cpu_sfence_valid),
        .frontend_io_ptw_pmp_1_cfg_a(frontend_io_ptw_pmp_1_cfg_a),
        .frontend_io_ptw_pmp_1_cfg_w(frontend_io_ptw_pmp_1_cfg_w),
        .frontend_io_ptw_pmp_2_cfg_a(frontend_io_ptw_pmp_2_cfg_a),
        .frontend_io_ptw_pmp_6_cfg_a(frontend_io_ptw_pmp_6_cfg_a),
        .frontend_io_ptw_pmp_7_cfg_a(frontend_io_ptw_pmp_7_cfg_a),
        .frontend_io_ptw_ptbr_mode(frontend_io_ptw_ptbr_mode),
        .frontend_io_ptw_status_prv(frontend_io_ptw_status_prv),
        .hitsVec_4(\tlb/hitsVec_4 ),
        .host_clk(host_clk),
        .ibuf_io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
        .ibuf_io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
        .ibuf_io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
        .ibuf_io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw[29]),
        .ibuf_io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
        .id_ctrl_fence_i(id_ctrl_fence_i),
        .id_ctrl_jal(id_ctrl_jal),
        .id_ctrl_mem(id_ctrl_mem),
        .id_ctrl_rxs2(id_ctrl_rxs2),
        .id_ctrl_sel_alu1(id_ctrl_sel_alu1),
        .id_ctrl_wxd(id_ctrl_wxd),
        .id_reg_fence_reg_0(core_n_1091),
        .invalidated(\icache/invalidated ),
        .invalidated_reg(core_n_680),
        .io_mask(fq_io_mask),
        .\lrscCount_reg[0] (core_n_1343),
        .\lrscCount_reg[0]_0 (core_n_1344),
        .mem_br_taken__reg_0(core_n_2317),
        .mem_ctrl_branch(mem_ctrl_branch),
        .mem_ctrl_branch_reg_0(core__710_n_0),
        .mem_ctrl_fence_i_reg_0(core__194_n_0),
        .mem_ctrl_fp(mem_ctrl_fp),
        .mem_ctrl_jal(mem_ctrl_jal),
        .mem_ctrl_jalr(mem_ctrl_jalr),
        .mem_ctrl_mem(mem_ctrl_mem),
        .mem_reg_flush_pipe(mem_reg_flush_pipe),
        .mem_reg_flush_pipe_reg_0(core__195_n_0),
        .\mem_reg_inst_reg[11]_0 (frontend_n_410),
        .\mem_reg_inst_reg[31]_0 ({_T_1686,core_n_1242,core_n_1243,dcacheArb_io_requestor_1_req_bits_tag}),
        .\mem_reg_inst_reg[9]_0 (core__691_n_0),
        .\mem_reg_inst_reg[9]_1 (ex_reg_rs_msb_0),
        .\mem_reg_pc_reg[31]_0 (ex_reg_pc),
        .mem_reg_replay_reg_0(mem_reg_replay_reg),
        .\mem_reg_rs2_reg[0]_0 (core_n_958),
        .\mem_reg_rs2_reg[1]_0 (core_n_959),
        .\mem_reg_rs2_reg[25]_0 (core_n_1775),
        .\mem_reg_rs2_reg[2]_0 (core_n_962),
        .\mem_reg_rs2_reg[3]_0 (core_n_964),
        .\mem_reg_rs2_reg[3]_1 ({core_n_1330,core_n_1331}),
        .\mem_reg_rs2_reg[4]_0 (core_n_965),
        .\mem_reg_rs2_reg[5]_0 (core_n_966),
        .\mem_reg_rs2_reg[6]_0 (core_n_906),
        .\mem_reg_rs2_reg[7]_0 (core_n_904),
        .mem_reg_rvc(mem_reg_rvc),
        .mem_reg_rvc_reg_0(core_n_16),
        .mem_reg_sfence(mem_reg_sfence),
        .mem_reg_sfence_reg_0(core_n_1364),
        .mem_reg_sfence_reg_1(core__193_n_0),
        .mem_reg_sfence_reg_2(core__201_n_0),
        .mem_reg_slow_bypass(mem_reg_slow_bypass),
        .mem_reg_slow_bypass_reg_0(core_n_1706),
        .mem_reg_slow_bypass_reg_1(core__196_n_0),
        .mem_reg_valid(mem_reg_valid),
        .mem_reg_valid_reg_0(core_n_1317),
        .mem_reg_xcpt(mem_reg_xcpt),
        .mem_reg_xcpt0(mem_reg_xcpt0),
        .mem_reg_xcpt_interrupt(mem_reg_xcpt_interrupt),
        .mem_reg_xcpt_interrupt_reg_0({core__709_n_0,core__708_n_0}),
        .nBufValid_reg(frontend_n_320),
        .nBufValid_reg_0(frontend_n_169),
        .nBufValid_reg_1(frontend_n_170),
        .nBufValid_reg_2(frontend_n_265),
        .nBufValid_reg_3(frontend_n_374),
        .nBufValid_reg_4(frontend_n_376),
        .nBufValid_reg_5(frontend_n_232),
        .nBufValid_reg_6(_T_1396__T_1405_addr),
        .nBufValid_reg_7(frontend_n_361),
        .nBufValid_reg_8(id_ctrl_sel_imm),
        .nBufValid_reg_9(\ibuf/_T_81 ),
        .neg_out_reg(core_n_289),
        .out({\trig_pc_reg[63]_i_2_n_4 ,\trig_pc_reg[63]_i_2_n_5 ,\trig_pc_reg[63]_i_2_n_6 ,\trig_pc_reg[63]_i_2_n_7 ,\trig_pc_reg[59]_i_1_n_4 ,\trig_pc_reg[59]_i_1_n_5 ,\trig_pc_reg[59]_i_1_n_6 ,\trig_pc_reg[59]_i_1_n_7 ,\trig_pc_reg[55]_i_1_n_4 ,\trig_pc_reg[55]_i_1_n_5 ,\trig_pc_reg[55]_i_1_n_6 ,\trig_pc_reg[55]_i_1_n_7 ,\trig_pc_reg[51]_i_1_n_4 ,\trig_pc_reg[51]_i_1_n_5 ,\trig_pc_reg[51]_i_1_n_6 ,\trig_pc_reg[51]_i_1_n_7 ,\trig_pc_reg[47]_i_1_n_4 ,\trig_pc_reg[47]_i_1_n_5 ,\trig_pc_reg[47]_i_1_n_6 ,\trig_pc_reg[47]_i_1_n_7 ,\trig_pc_reg[43]_i_1_n_4 ,\trig_pc_reg[43]_i_1_n_5 ,\trig_pc_reg[43]_i_1_n_6 ,\trig_pc_reg[43]_i_1_n_7 ,\trig_pc_reg[39]_i_1_n_4 ,\trig_pc_reg[39]_i_1_n_5 ,\trig_pc_reg[39]_i_1_n_6 ,\trig_pc_reg[39]_i_1_n_7 ,\trig_pc_reg[35]_i_1_n_4 ,\trig_pc_reg[35]_i_1_n_5 ,\trig_pc_reg[35]_i_1_n_6 ,\trig_pc_reg[35]_i_1_n_7 ,\trig_pc_reg[31]_i_1_n_4 ,\trig_pc_reg[31]_i_1_n_5 ,\trig_pc_reg[31]_i_1_n_6 ,\trig_pc_reg[31]_i_1_n_7 ,\trig_pc_reg[27]_i_1_n_4 ,\trig_pc_reg[27]_i_1_n_5 ,\trig_pc_reg[27]_i_1_n_6 ,\trig_pc_reg[27]_i_1_n_7 ,\trig_pc_reg[23]_i_1_n_4 ,\trig_pc_reg[23]_i_1_n_5 ,\trig_pc_reg[23]_i_1_n_6 ,\trig_pc_reg[23]_i_1_n_7 ,\trig_pc_reg[19]_i_1_n_4 ,\trig_pc_reg[19]_i_1_n_5 ,\trig_pc_reg[19]_i_1_n_6 ,\trig_pc_reg[19]_i_1_n_7 ,\trig_pc_reg[15]_i_1_n_4 ,\trig_pc_reg[15]_i_1_n_5 ,\trig_pc_reg[15]_i_1_n_6 ,\trig_pc_reg[15]_i_1_n_7 ,\trig_pc_reg[11]_i_1_n_4 ,\trig_pc_reg[11]_i_1_n_5 ,\trig_pc_reg[11]_i_1_n_6 ,\trig_pc_reg[11]_i_1_n_7 ,\trig_pc_reg[7]_i_1_n_4 ,\trig_pc_reg[7]_i_1_n_5 ,\trig_pc_reg[7]_i_1_n_6 ,\trig_pc_reg[7]_i_1_n_7 ,\trig_pc_reg[3]_i_1_n_4 ,\trig_pc_reg[3]_i_1_n_5 ,\trig_pc_reg[3]_i_1_n_6 ,\trig_pc_reg[3]_i_1_n_7 }),
        .p_0_in(p_0_in),
        .p_13_in(\tlb/p_13_in ),
        .p_2_in(\tlb/p_2_in ),
        .p_31_in(p_31_in),
        .q_reg(q_reg),
        .\r_pte_ppn_reg[0] (ptw_n_15),
        .\r_pte_ppn_reg[10] (ptw_n_183),
        .\r_pte_ppn_reg[11] (ptw_n_162),
        .\r_pte_ppn_reg[12] (ptw_n_170),
        .\r_pte_ppn_reg[13] (ptw_n_167),
        .\r_pte_ppn_reg[14] (ptw_n_168),
        .\r_pte_ppn_reg[15] (ptw_n_160),
        .\r_pte_ppn_reg[16] (ptw_n_89),
        .\r_pte_ppn_reg[16]_0 (ptw_n_94),
        .\r_pte_ppn_reg[16]_1 (ptw_n_98),
        .\r_pte_ppn_reg[16]_2 (ptw_n_102),
        .\r_pte_ppn_reg[16]_3 (ptw_n_107),
        .\r_pte_ppn_reg[16]_4 (ptw_n_112),
        .\r_pte_ppn_reg[16]_5 (ptw_n_117),
        .\r_pte_ppn_reg[16]_6 (ptw_n_122),
        .\r_pte_ppn_reg[16]_7 (ptw_n_161),
        .\r_pte_ppn_reg[17] (ptw_n_163),
        .\r_pte_ppn_reg[18] (ptw_n_134),
        .\r_pte_ppn_reg[19] (ptw_io_dpath_ptbr_ppn),
        .\r_pte_ppn_reg[19]_0 (dcache_io_ptw_resp_bits_pte_ppn),
        .\r_pte_ppn_reg[1] (ptw_n_14),
        .\r_pte_ppn_reg[2] (ptw_n_13),
        .\r_pte_ppn_reg[3] (ptw_n_86),
        .\r_pte_ppn_reg[3]_0 (ptw_n_91),
        .\r_pte_ppn_reg[3]_1 (ptw_n_95),
        .\r_pte_ppn_reg[3]_2 (ptw_n_99),
        .\r_pte_ppn_reg[3]_3 (ptw_n_104),
        .\r_pte_ppn_reg[3]_4 (ptw_n_109),
        .\r_pte_ppn_reg[3]_5 (ptw_n_114),
        .\r_pte_ppn_reg[3]_6 (ptw_n_119),
        .\r_pte_ppn_reg[3]_7 (ptw_n_173),
        .\r_pte_ppn_reg[4] (ptw_n_172),
        .\r_pte_ppn_reg[5] (ptw_n_174),
        .\r_pte_ppn_reg[5]_0 (ptw_n_87),
        .\r_pte_ppn_reg[5]_1 (ptw_n_92),
        .\r_pte_ppn_reg[5]_2 (ptw_n_96),
        .\r_pte_ppn_reg[5]_3 (ptw_n_100),
        .\r_pte_ppn_reg[5]_4 (ptw_n_105),
        .\r_pte_ppn_reg[5]_5 (ptw_n_110),
        .\r_pte_ppn_reg[5]_6 (ptw_n_115),
        .\r_pte_ppn_reg[5]_7 (ptw_n_120),
        .\r_pte_ppn_reg[6] (ptw_n_176),
        .\r_pte_ppn_reg[7] (ptw_n_88),
        .\r_pte_ppn_reg[7]_0 (ptw_n_93),
        .\r_pte_ppn_reg[7]_1 (ptw_n_97),
        .\r_pte_ppn_reg[7]_2 (ptw_n_101),
        .\r_pte_ppn_reg[7]_3 (ptw_n_106),
        .\r_pte_ppn_reg[7]_4 (ptw_n_111),
        .\r_pte_ppn_reg[7]_5 (ptw_n_116),
        .\r_pte_ppn_reg[7]_6 (ptw_n_121),
        .\r_pte_ppn_reg[7]_7 (ptw_n_178),
        .\r_pte_ppn_reg[8] (ptw_n_177),
        .\r_pte_ppn_reg[9] (ptw_n_182),
        .\r_refill_waddr_reg[0] (core_n_1840),
        .\r_refill_waddr_reg[1] ({frontend_n_51,frontend_n_52}),
        .refill_valid(\icache/refill_valid ),
        .\reg_bp_0_address_reg[36] (\bpu/_T_132 ),
        .\reg_bp_0_address_reg[3] (core__127_n_0),
        .reg_bp_0_control_action_reg(core__128_n_0),
        .\reg_bp_0_control_tmatch_reg[1] ({csr_io_rw_addr[11:9],csr_io_rw_addr[7:6],csr_io_rw_addr[4],csr_io_rw_addr[2:0],wb_waddr}),
        .\reg_bp_0_control_tmatch_reg[1]_0 (core_n_1018),
        .\reg_dcsr_cause_reg[0] (core_n_1014),
        .\reg_dcsr_cause_reg[1] (core_n_1009),
        .reg_dcsr_prv(\csr/reg_dcsr_prv ),
        .reg_dcsr_step(\csr/reg_dcsr_step ),
        .reg_debug_reg(core_n_1003),
        .reg_debug_reg_0(core__107_n_0),
        .reg_debug_reg_1(core__102_n_0),
        .reg_debug_reg_2(core__120_n_0),
        .\reg_dpc_reg[12] (core_n_947),
        .\reg_dpc_reg[39] (wb_reg_pc),
        .\reg_dscratch_reg[0] (core_n_957),
        .\reg_entries_0_reg[0] (core_n_423),
        .\reg_entries_0_reg[0]_0 (core_n_809),
        .\reg_entries_0_reg[0]_1 (core_n_883),
        .\reg_entries_0_reg[0]_2 (core_n_884),
        .\reg_entries_0_reg[0]_3 (core_n_885),
        .\reg_entries_0_reg[0]_4 (core_n_886),
        .\reg_entries_0_reg[0]_5 (core_n_887),
        .\reg_entries_0_reg[0]_6 (core_n_888),
        .\reg_entries_0_reg[0]_7 (core_n_889),
        .\reg_entries_0_reg[10] (\tlb/_GEN_36 ),
        .\reg_entries_0_reg[4] (core_n_1835),
        .\reg_entries_0_reg[4]_0 (core_n_1843),
        .\reg_entries_0_reg[4]_1 ({core_n_1844,core_n_1845,core_n_1846}),
        .\reg_entries_0_reg[4]_10 ({core_n_1971,core_n_1972,core_n_1973,core_n_1974}),
        .\reg_entries_0_reg[4]_11 ({core_n_1975,core_n_1976,core_n_1977,core_n_1978}),
        .\reg_entries_0_reg[4]_12 ({core_n_1979,core_n_1980,core_n_1981,core_n_1982}),
        .\reg_entries_0_reg[4]_13 ({core_n_1994,core_n_1995,core_n_1996}),
        .\reg_entries_0_reg[4]_14 (core_n_2003),
        .\reg_entries_0_reg[4]_15 (core_n_2004),
        .\reg_entries_0_reg[4]_16 (core_n_2005),
        .\reg_entries_0_reg[4]_17 (core_n_2033),
        .\reg_entries_0_reg[4]_18 (core_n_2051),
        .\reg_entries_0_reg[4]_19 (core_n_2060),
        .\reg_entries_0_reg[4]_2 ({core_n_1847,core_n_1848,core_n_1849}),
        .\reg_entries_0_reg[4]_20 ({core_n_2061,core_n_2062,core_n_2063,core_n_2064}),
        .\reg_entries_0_reg[4]_21 ({core_n_2065,core_n_2066,core_n_2067,core_n_2068}),
        .\reg_entries_0_reg[4]_22 (core_n_2069),
        .\reg_entries_0_reg[4]_23 ({core_n_2070,core_n_2071,core_n_2072,core_n_2073}),
        .\reg_entries_0_reg[4]_24 ({core_n_2074,core_n_2075,core_n_2076,core_n_2077}),
        .\reg_entries_0_reg[4]_25 (core_n_2078),
        .\reg_entries_0_reg[4]_3 ({core_n_1875,core_n_1876}),
        .\reg_entries_0_reg[4]_4 ({core_n_1877,core_n_1878}),
        .\reg_entries_0_reg[4]_5 ({core_n_1915,core_n_1916,core_n_1917,core_n_1918}),
        .\reg_entries_0_reg[4]_6 ({core_n_1919,core_n_1920,core_n_1921,core_n_1922}),
        .\reg_entries_0_reg[4]_7 ({core_n_1923,core_n_1924,core_n_1925,core_n_1926}),
        .\reg_entries_0_reg[4]_8 (core_n_1927),
        .\reg_entries_0_reg[4]_9 ({core_n_1928,core_n_1929,core_n_1930,core_n_1931}),
        .\reg_entries_0_reg[5] (\tlb/_T_952 ),
        .\reg_entries_0_reg[5]_0 ({core_n_692,core_n_693,core_n_694,core_n_695}),
        .\reg_entries_0_reg[5]_1 ({core_n_700,core_n_701,core_n_702,core_n_703}),
        .\reg_entries_0_reg[5]_10 ({core_n_759,core_n_760,core_n_761}),
        .\reg_entries_0_reg[5]_11 ({core_n_762,core_n_763,core_n_764}),
        .\reg_entries_0_reg[5]_12 ({core_n_765,core_n_766,core_n_767}),
        .\reg_entries_0_reg[5]_13 ({core_n_768,core_n_769,core_n_770}),
        .\reg_entries_0_reg[5]_14 ({core_n_771,core_n_772,core_n_773}),
        .\reg_entries_0_reg[5]_15 ({core_n_774,core_n_775,core_n_776}),
        .\reg_entries_0_reg[5]_16 ({core_n_777,core_n_778,core_n_779,core_n_780}),
        .\reg_entries_0_reg[5]_17 ({core_n_781,core_n_782,core_n_783,core_n_784}),
        .\reg_entries_0_reg[5]_18 ({core_n_785,core_n_786,core_n_787,core_n_788}),
        .\reg_entries_0_reg[5]_19 ({core_n_789,core_n_790,core_n_791,core_n_792}),
        .\reg_entries_0_reg[5]_2 ({core_n_708,core_n_709,core_n_710,core_n_711}),
        .\reg_entries_0_reg[5]_20 ({core_n_793,core_n_794,core_n_795,core_n_796}),
        .\reg_entries_0_reg[5]_21 ({core_n_797,core_n_798,core_n_799,core_n_800}),
        .\reg_entries_0_reg[5]_22 ({core_n_801,core_n_802,core_n_803,core_n_804}),
        .\reg_entries_0_reg[5]_23 ({core_n_805,core_n_806,core_n_807,core_n_808}),
        .\reg_entries_0_reg[5]_24 ({core_n_811,core_n_812,core_n_813,core_n_814}),
        .\reg_entries_0_reg[5]_25 ({core_n_815,core_n_816,core_n_817,core_n_818}),
        .\reg_entries_0_reg[5]_26 (core_n_819),
        .\reg_entries_0_reg[5]_27 ({core_n_820,core_n_821,core_n_822,core_n_823}),
        .\reg_entries_0_reg[5]_28 ({core_n_824,core_n_825,core_n_826,core_n_827}),
        .\reg_entries_0_reg[5]_29 (core_n_828),
        .\reg_entries_0_reg[5]_3 ({core_n_712,core_n_713,core_n_714,core_n_715}),
        .\reg_entries_0_reg[5]_30 ({core_n_829,core_n_830,core_n_831,core_n_832}),
        .\reg_entries_0_reg[5]_31 ({core_n_833,core_n_834,core_n_835,core_n_836}),
        .\reg_entries_0_reg[5]_32 (core_n_837),
        .\reg_entries_0_reg[5]_33 ({core_n_838,core_n_839,core_n_840,core_n_841}),
        .\reg_entries_0_reg[5]_34 ({core_n_842,core_n_843,core_n_844,core_n_845}),
        .\reg_entries_0_reg[5]_35 (core_n_846),
        .\reg_entries_0_reg[5]_36 ({core_n_847,core_n_848,core_n_849,core_n_850}),
        .\reg_entries_0_reg[5]_37 ({core_n_851,core_n_852,core_n_853,core_n_854}),
        .\reg_entries_0_reg[5]_38 (core_n_855),
        .\reg_entries_0_reg[5]_39 ({core_n_856,core_n_857,core_n_858,core_n_859}),
        .\reg_entries_0_reg[5]_4 ({core_n_721,core_n_722,core_n_723,core_n_724}),
        .\reg_entries_0_reg[5]_40 ({core_n_860,core_n_861,core_n_862,core_n_863}),
        .\reg_entries_0_reg[5]_41 (core_n_864),
        .\reg_entries_0_reg[5]_42 ({core_n_865,core_n_866,core_n_867,core_n_868}),
        .\reg_entries_0_reg[5]_43 ({core_n_869,core_n_870,core_n_871,core_n_872}),
        .\reg_entries_0_reg[5]_44 (core_n_873),
        .\reg_entries_0_reg[5]_45 ({core_n_874,core_n_875,core_n_876,core_n_877}),
        .\reg_entries_0_reg[5]_46 ({core_n_878,core_n_879,core_n_880,core_n_881}),
        .\reg_entries_0_reg[5]_47 (core_n_882),
        .\reg_entries_0_reg[5]_5 ({core_n_730,core_n_731,core_n_732,core_n_733}),
        .\reg_entries_0_reg[5]_6 ({core_n_736,core_n_737,core_n_738,core_n_739}),
        .\reg_entries_0_reg[5]_7 ({core_n_745,core_n_746,core_n_747,core_n_748}),
        .\reg_entries_0_reg[5]_8 ({core_n_753,core_n_754,core_n_755}),
        .\reg_entries_0_reg[5]_9 ({core_n_756,core_n_757,core_n_758}),
        .\reg_entries_0_reg[6] ({core_n_391,core_n_392,core_n_393}),
        .\reg_entries_0_reg[6]_0 ({core_n_424,core_n_425,core_n_426}),
        .\reg_entries_0_reg[6]_1 (core_n_459),
        .\reg_entries_0_reg[6]_10 ({core_n_1856,core_n_1857,core_n_1858}),
        .\reg_entries_0_reg[6]_11 ({core_n_1859,core_n_1860,core_n_1861}),
        .\reg_entries_0_reg[6]_12 ({core_n_1862,core_n_1863,core_n_1864}),
        .\reg_entries_0_reg[6]_13 ({core_n_1865,core_n_1866,core_n_1867}),
        .\reg_entries_0_reg[6]_14 (core_n_1868),
        .\reg_entries_0_reg[6]_15 ({core_n_1869,core_n_1870}),
        .\reg_entries_0_reg[6]_16 ({core_n_1871,core_n_1872}),
        .\reg_entries_0_reg[6]_17 ({core_n_1873,core_n_1874}),
        .\reg_entries_0_reg[6]_18 ({core_n_1879,core_n_1880,core_n_1881,core_n_1882}),
        .\reg_entries_0_reg[6]_19 ({core_n_1883,core_n_1884,core_n_1885,core_n_1886}),
        .\reg_entries_0_reg[6]_2 (core_n_518),
        .\reg_entries_0_reg[6]_20 ({core_n_1887,core_n_1888,core_n_1889,core_n_1890}),
        .\reg_entries_0_reg[6]_21 ({core_n_1891,core_n_1892,core_n_1893,core_n_1894}),
        .\reg_entries_0_reg[6]_22 ({core_n_1895,core_n_1896,core_n_1897,core_n_1898}),
        .\reg_entries_0_reg[6]_23 ({core_n_1899,core_n_1900,core_n_1901,core_n_1902}),
        .\reg_entries_0_reg[6]_24 ({core_n_1903,core_n_1904,core_n_1905,core_n_1906}),
        .\reg_entries_0_reg[6]_25 ({core_n_1907,core_n_1908,core_n_1909,core_n_1910}),
        .\reg_entries_0_reg[6]_26 ({core_n_1911,core_n_1912,core_n_1913,core_n_1914}),
        .\reg_entries_0_reg[6]_27 ({core_n_1932,core_n_1933,core_n_1934}),
        .\reg_entries_0_reg[6]_28 ({core_n_1935,core_n_1936,core_n_1937,core_n_1938}),
        .\reg_entries_0_reg[6]_29 ({core_n_1939,core_n_1940,core_n_1941,core_n_1942}),
        .\reg_entries_0_reg[6]_3 (core_n_519),
        .\reg_entries_0_reg[6]_30 ({core_n_1943,core_n_1944,core_n_1945,core_n_1946}),
        .\reg_entries_0_reg[6]_31 ({core_n_1947,core_n_1948,core_n_1949,core_n_1950}),
        .\reg_entries_0_reg[6]_32 ({core_n_1951,core_n_1952,core_n_1953,core_n_1954}),
        .\reg_entries_0_reg[6]_33 ({core_n_1955,core_n_1956,core_n_1957,core_n_1958}),
        .\reg_entries_0_reg[6]_34 ({core_n_1959,core_n_1960,core_n_1961,core_n_1962}),
        .\reg_entries_0_reg[6]_35 ({core_n_1963,core_n_1964,core_n_1965,core_n_1966}),
        .\reg_entries_0_reg[6]_36 ({core_n_1967,core_n_1968,core_n_1969,core_n_1970}),
        .\reg_entries_0_reg[6]_37 ({core_n_1983,core_n_1984,core_n_1985,core_n_1986}),
        .\reg_entries_0_reg[6]_38 ({core_n_1987,core_n_1988,core_n_1989}),
        .\reg_entries_0_reg[6]_39 ({core_n_1990,core_n_1991,core_n_1992,core_n_1993}),
        .\reg_entries_0_reg[6]_4 (core_n_520),
        .\reg_entries_0_reg[6]_40 ({core_n_1997,core_n_1998,core_n_1999}),
        .\reg_entries_0_reg[6]_41 ({core_n_2000,core_n_2001,core_n_2002}),
        .\reg_entries_0_reg[6]_42 (core_n_2006),
        .\reg_entries_0_reg[6]_43 ({core_n_2007,core_n_2008,core_n_2009,core_n_2010}),
        .\reg_entries_0_reg[6]_44 ({core_n_2011,core_n_2012,core_n_2013,core_n_2014}),
        .\reg_entries_0_reg[6]_45 (core_n_2015),
        .\reg_entries_0_reg[6]_46 ({core_n_2016,core_n_2017,core_n_2018,core_n_2019}),
        .\reg_entries_0_reg[6]_47 ({core_n_2020,core_n_2021,core_n_2022,core_n_2023}),
        .\reg_entries_0_reg[6]_48 (core_n_2024),
        .\reg_entries_0_reg[6]_49 ({core_n_2025,core_n_2026,core_n_2027,core_n_2028}),
        .\reg_entries_0_reg[6]_5 ({\tlb/_T_949 ,\tlb/_T_946 }),
        .\reg_entries_0_reg[6]_50 ({core_n_2029,core_n_2030,core_n_2031,core_n_2032}),
        .\reg_entries_0_reg[6]_51 ({core_n_2034,core_n_2035,core_n_2036,core_n_2037}),
        .\reg_entries_0_reg[6]_52 ({core_n_2038,core_n_2039,core_n_2040,core_n_2041}),
        .\reg_entries_0_reg[6]_53 (core_n_2042),
        .\reg_entries_0_reg[6]_54 ({core_n_2043,core_n_2044,core_n_2045,core_n_2046}),
        .\reg_entries_0_reg[6]_55 ({core_n_2047,core_n_2048,core_n_2049,core_n_2050}),
        .\reg_entries_0_reg[6]_56 ({core_n_2052,core_n_2053,core_n_2054,core_n_2055}),
        .\reg_entries_0_reg[6]_57 ({core_n_2056,core_n_2057,core_n_2058,core_n_2059}),
        .\reg_entries_0_reg[6]_6 (core_n_1836),
        .\reg_entries_0_reg[6]_7 (core_n_1842),
        .\reg_entries_0_reg[6]_8 ({core_n_1850,core_n_1851,core_n_1852}),
        .\reg_entries_0_reg[6]_9 ({core_n_1853,core_n_1854,core_n_1855}),
        .\reg_entries_1_reg[0] (core_n_639),
        .\reg_entries_1_reg[0]_0 (core_n_640),
        .\reg_entries_1_reg[0]_1 (core_n_641),
        .\reg_entries_1_reg[0]_10 ({frontend_io_ptw_pmp_5_mask[29],frontend_io_ptw_pmp_5_mask[20],frontend_io_ptw_pmp_5_mask[11]}),
        .\reg_entries_1_reg[0]_11 ({frontend_io_ptw_pmp_4_mask[29],frontend_io_ptw_pmp_4_mask[20],frontend_io_ptw_pmp_4_mask[11]}),
        .\reg_entries_1_reg[0]_12 ({frontend_io_ptw_pmp_7_mask[29],frontend_io_ptw_pmp_7_mask[20],frontend_io_ptw_pmp_7_mask[11]}),
        .\reg_entries_1_reg[0]_13 ({frontend_io_ptw_pmp_6_mask[29],frontend_io_ptw_pmp_6_mask[20],frontend_io_ptw_pmp_6_mask[11]}),
        .\reg_entries_1_reg[0]_14 ({frontend_io_ptw_pmp_1_mask[29],frontend_io_ptw_pmp_1_mask[20],frontend_io_ptw_pmp_1_mask[11]}),
        .\reg_entries_1_reg[0]_15 (core_n_1800),
        .\reg_entries_1_reg[0]_16 (core_n_1801),
        .\reg_entries_1_reg[0]_17 (core_n_1802),
        .\reg_entries_1_reg[0]_18 (core_n_1803),
        .\reg_entries_1_reg[0]_19 (core_n_1804),
        .\reg_entries_1_reg[0]_2 (core_n_642),
        .\reg_entries_1_reg[0]_20 (core_n_1805),
        .\reg_entries_1_reg[0]_21 (core_n_1806),
        .\reg_entries_1_reg[0]_22 (core_n_1807),
        .\reg_entries_1_reg[0]_23 (core_n_1808),
        .\reg_entries_1_reg[0]_24 (core_n_1809),
        .\reg_entries_1_reg[0]_25 (core_n_1810),
        .\reg_entries_1_reg[0]_26 (core_n_1811),
        .\reg_entries_1_reg[0]_27 (core_n_1812),
        .\reg_entries_1_reg[0]_28 (core_n_1813),
        .\reg_entries_1_reg[0]_29 (core_n_1814),
        .\reg_entries_1_reg[0]_3 (core_n_643),
        .\reg_entries_1_reg[0]_30 (core_n_1815),
        .\reg_entries_1_reg[0]_31 (core_n_1816),
        .\reg_entries_1_reg[0]_32 (core_n_1817),
        .\reg_entries_1_reg[0]_33 (core_n_1818),
        .\reg_entries_1_reg[0]_34 (core_n_1819),
        .\reg_entries_1_reg[0]_35 (core_n_1820),
        .\reg_entries_1_reg[0]_36 (core_n_1821),
        .\reg_entries_1_reg[0]_37 (core_n_1822),
        .\reg_entries_1_reg[0]_38 (core_n_1823),
        .\reg_entries_1_reg[0]_39 (core_n_1824),
        .\reg_entries_1_reg[0]_4 (core_n_644),
        .\reg_entries_1_reg[0]_40 (core_n_1825),
        .\reg_entries_1_reg[0]_41 (core_n_1826),
        .\reg_entries_1_reg[0]_42 (core_n_1827),
        .\reg_entries_1_reg[0]_43 (core_n_1828),
        .\reg_entries_1_reg[0]_44 (core_n_1829),
        .\reg_entries_1_reg[0]_45 (core_n_1830),
        .\reg_entries_1_reg[0]_46 (core_n_1831),
        .\reg_entries_1_reg[0]_47 (core_n_1832),
        .\reg_entries_1_reg[0]_5 (core_n_645),
        .\reg_entries_1_reg[0]_6 (core_n_646),
        .\reg_entries_1_reg[0]_7 (core_n_649),
        .\reg_entries_1_reg[0]_8 ({frontend_io_ptw_pmp_2_mask[29],frontend_io_ptw_pmp_2_mask[20],frontend_io_ptw_pmp_2_mask[11]}),
        .\reg_entries_1_reg[0]_9 (core_n_687),
        .\reg_entries_1_reg[12] (\tlb/entries_1_u ),
        .\reg_entries_2_reg[12] ({\tlb/entries_2_u ,\tlb/entries_2_sx ,\tlb/entries_2_sr }),
        .\reg_entries_3_reg[11] (\tlb/entries_3_g ),
        .\reg_entries_3_reg[12] ({\tlb/entries_3_u ,\tlb/entries_3_sx ,\tlb/entries_3_sr }),
        .\reg_entries_4_reg[61] ({\tlb/p_0_in [19:18],\tlb/p_0_in [14],\tlb/p_0_in [12],\tlb/p_0_in [8],\tlb/p_0_in [6],\tlb/p_0_in [0],\tlb/entries_4_u ,\tlb/entries_4_sx ,\tlb/entries_4_sr }),
        .\reg_entries_4_reg[61]_0 (dcache_n_585),
        .\reg_mbadaddr_reg[12] (core_n_902),
        .\reg_mcause_reg[0] (core_n_963),
        .\reg_mepc_reg[12] (core_n_909),
        .\reg_mie_reg[7] (Q),
        .reg_mip_seip_reg(core_n_895),
        .reg_mip_seip_reg_0(core_n_910),
        .\reg_misa_reg[0] (core_n_994),
        .\reg_misa_reg[12] ({csr_io_status_isa[12],csr_io_status_isa[2]}),
        .\reg_misa_reg[12]_0 (frontend_n_356),
        .reg_mstatus_mie(\csr/reg_mstatus_mie ),
        .reg_mstatus_mie_reg(core_n_999),
        .reg_mstatus_mie_reg_0(core_n_1008),
        .reg_mstatus_mpie_reg(core_n_86),
        .reg_mstatus_mpie_reg_0(core_n_1005),
        .\reg_mstatus_mpp_reg[0] (core_n_1007),
        .\reg_mstatus_mpp_reg[1] (core_n_1006),
        .\reg_mstatus_prv_reg[1] (core_n_1004),
        .\reg_mstatus_prv_reg[1]_0 (core__117_n_0),
        .\reg_mstatus_prv_reg[1]_1 (core__126_n_0),
        .\reg_mstatus_prv_reg[1]_2 (core__129_n_0),
        .reg_mstatus_spie_reg(core_n_85),
        .reg_mstatus_tvm_reg(frontend_n_352),
        .\reg_mtvec_reg[10] (core_n_912),
        .\reg_mtvec_reg[11] (core_n_913),
        .\reg_mtvec_reg[12] (core_n_897),
        .\reg_mtvec_reg[13] (core_n_914),
        .\reg_mtvec_reg[14] (core_n_940),
        .\reg_mtvec_reg[15] (core_n_941),
        .\reg_mtvec_reg[16] (core_n_942),
        .\reg_mtvec_reg[17] (core_n_943),
        .\reg_mtvec_reg[18] (core_n_944),
        .\reg_mtvec_reg[19] (core_n_945),
        .\reg_mtvec_reg[20] (core_n_68),
        .\reg_mtvec_reg[20]_0 (core_n_946),
        .\reg_mtvec_reg[21] (core_n_69),
        .\reg_mtvec_reg[21]_0 (core_n_948),
        .\reg_mtvec_reg[22] (core_n_70),
        .\reg_mtvec_reg[22]_0 (core_n_949),
        .\reg_mtvec_reg[23] (core_n_950),
        .\reg_mtvec_reg[24] (core_n_951),
        .\reg_mtvec_reg[25] (core_n_952),
        .\reg_mtvec_reg[26] (core_n_953),
        .\reg_mtvec_reg[27] (core_n_954),
        .\reg_mtvec_reg[28] (core_n_955),
        .\reg_mtvec_reg[29] ({frontend_io_ptw_pmp_1_addr[29:7],frontend_io_ptw_pmp_1_addr[5:0]}),
        .\reg_mtvec_reg[29]_0 (frontend_io_ptw_pmp_2_addr),
        .\reg_mtvec_reg[29]_1 ({frontend_io_ptw_pmp_3_addr[29:10],frontend_io_ptw_pmp_3_addr[8:7],frontend_io_ptw_pmp_3_addr[5:0]}),
        .\reg_mtvec_reg[29]_2 (frontend_io_ptw_pmp_0_addr),
        .\reg_mtvec_reg[29]_3 (frontend_io_ptw_pmp_4_addr),
        .\reg_mtvec_reg[29]_4 ({frontend_io_ptw_pmp_7_addr[29:10],frontend_io_ptw_pmp_7_addr[8:7],frontend_io_ptw_pmp_7_addr[5:0]}),
        .\reg_mtvec_reg[29]_5 ({frontend_io_ptw_pmp_6_addr[29:3],frontend_io_ptw_pmp_6_addr[1:0]}),
        .\reg_mtvec_reg[29]_6 ({frontend_io_ptw_pmp_5_addr[29:5],frontend_io_ptw_pmp_5_addr[3:0]}),
        .\reg_mtvec_reg[29]_7 (core_n_956),
        .\reg_mtvec_reg[30] (core_n_976),
        .\reg_mtvec_reg[31] (core_n_975),
        .\reg_mtvec_reg[4] (core__116_n_0),
        .\reg_mtvec_reg[8] (core_n_908),
        .\reg_pmp_0_addr_reg[13] (frontend_n_151),
        .\reg_pmp_0_addr_reg[17] (frontend_n_134),
        .\reg_pmp_0_addr_reg[19] (frontend_n_143),
        .\reg_pmp_0_addr_reg[23] (ptw_n_153),
        .\reg_pmp_0_addr_reg[28] (\tlb/pmp/_T_269 ),
        .\reg_pmp_0_addr_reg[28]_0 (_T_963),
        .\reg_pmp_0_addr_reg[29] (frontend_n_114),
        .\reg_pmp_0_addr_reg[29]_0 (\tlb/pmp/_T_836 ),
        .\reg_pmp_1_addr_reg[13] (frontend_n_150),
        .\reg_pmp_1_addr_reg[17] (frontend_n_133),
        .\reg_pmp_1_addr_reg[19] (frontend_n_142),
        .\reg_pmp_1_addr_reg[28] (\tlb/pmp/_T_233 ),
        .\reg_pmp_1_addr_reg[28]_0 (_T_1038),
        .\reg_pmp_1_addr_reg[29] (frontend_n_115),
        .\reg_pmp_1_addr_reg[29]_0 (\tlb/pmp/_T_709 ),
        .\reg_pmp_1_cfg_a_reg[0] (dcache_n_614),
        .reg_pmp_1_cfg_w_reg(dcache_n_613),
        .\reg_pmp_2_addr_reg[0] (ptw_n_139),
        .\reg_pmp_2_addr_reg[13] (frontend_n_149),
        .\reg_pmp_2_addr_reg[17] (frontend_n_132),
        .\reg_pmp_2_addr_reg[19] (frontend_n_141),
        .\reg_pmp_2_addr_reg[28] (\tlb/pmp/_T_197 ),
        .\reg_pmp_2_addr_reg[28]_0 (_T_1113),
        .\reg_pmp_2_addr_reg[29] (core_n_996),
        .\reg_pmp_2_addr_reg[29]_0 (frontend_n_116),
        .\reg_pmp_2_addr_reg[29]_1 (\tlb/pmp/_T_582 ),
        .\reg_pmp_2_cfg_a_reg[0] (dcache_n_616),
        .\reg_pmp_3_addr_reg[13] (frontend_n_146),
        .\reg_pmp_3_addr_reg[17] (frontend_n_129),
        .\reg_pmp_3_addr_reg[18] (ptw_n_181),
        .\reg_pmp_3_addr_reg[19] (frontend_n_138),
        .\reg_pmp_3_addr_reg[23] (ptw_n_169),
        .\reg_pmp_3_addr_reg[28] (\tlb/pmp/_T_161 ),
        .\reg_pmp_3_addr_reg[28]_0 (_T_1188),
        .\reg_pmp_3_addr_reg[29] (frontend_n_119),
        .\reg_pmp_3_addr_reg[29]_0 (\tlb/pmp/_T_455 ),
        .\reg_pmp_3_addr_reg[29]_1 (ptw_n_146),
        .\reg_pmp_4_addr_reg[0] (ptw_n_142),
        .\reg_pmp_4_addr_reg[13] (frontend_n_145),
        .\reg_pmp_4_addr_reg[14] (ptw_n_143),
        .\reg_pmp_4_addr_reg[17] (frontend_n_128),
        .\reg_pmp_4_addr_reg[19] (frontend_n_137),
        .\reg_pmp_4_addr_reg[28] (\tlb/pmp/_T_125 ),
        .\reg_pmp_4_addr_reg[28]_0 (_T_1263),
        .\reg_pmp_4_addr_reg[29] (frontend_n_120),
        .\reg_pmp_4_addr_reg[29]_0 (\tlb/pmp/_T_328 ),
        .\reg_pmp_4_cfg_a_reg[1] (frontend_io_ptw_pmp_4_cfg_a),
        .\reg_pmp_5_addr_reg[13] (frontend_n_144),
        .\reg_pmp_5_addr_reg[17] (frontend_n_127),
        .\reg_pmp_5_addr_reg[19] (frontend_n_136),
        .\reg_pmp_5_addr_reg[20] (core__111_n_0),
        .\reg_pmp_5_addr_reg[28] (\tlb/pmp/_T_89 ),
        .\reg_pmp_5_addr_reg[28]_0 (_T_1338),
        .\reg_pmp_5_addr_reg[29] (frontend_n_121),
        .\reg_pmp_5_addr_reg[29]_0 (\tlb/pmp/_T_201 ),
        .\reg_pmp_5_cfg_a_reg[1] (frontend_io_ptw_pmp_5_cfg_a),
        .\reg_pmp_5_cfg_a_reg[1]_0 (ptw_n_77),
        .\reg_pmp_6_addr_reg[13] (frontend_n_148),
        .\reg_pmp_6_addr_reg[17] (frontend_n_131),
        .\reg_pmp_6_addr_reg[19] (frontend_n_140),
        .\reg_pmp_6_addr_reg[28] (\tlb/pmp/_T_53 ),
        .\reg_pmp_6_addr_reg[28]_0 (_T_1413),
        .\reg_pmp_6_addr_reg[29] (frontend_n_117),
        .\reg_pmp_6_addr_reg[29]_0 (\tlb/pmp/_T_74 ),
        .\reg_pmp_7_addr_reg[13] (frontend_n_147),
        .\reg_pmp_7_addr_reg[17] (frontend_n_130),
        .\reg_pmp_7_addr_reg[17]_0 (ptw_n_180),
        .\reg_pmp_7_addr_reg[19] (frontend_n_139),
        .\reg_pmp_7_addr_reg[23] (ptw_n_171),
        .\reg_pmp_7_addr_reg[28] (\tlb/pmp/_T_58 ),
        .\reg_pmp_7_addr_reg[28]_0 (_T_1488),
        .\reg_pmp_7_addr_reg[29] (core_n_896),
        .\reg_pmp_7_addr_reg[29]_0 (frontend_n_118),
        .\reg_pmp_7_addr_reg[29]_1 (\tlb/pmp/_T_94 ),
        .\reg_pmp_7_addr_reg[29]_2 (ptw_n_159),
        .\reg_pmp_7_cfg_a_reg[0] (dcache_n_623),
        .\reg_sbadaddr_reg[0] (core_n_992),
        .\reg_sbadaddr_reg[30] ({core_n_1332,core_n_1333,core_n_1334}),
        .\reg_sbadaddr_reg[30]_0 ({core_n_1335,core_n_1336,core_n_1337}),
        .\reg_sbadaddr_reg[30]_1 ({core_n_1338,core_n_1339,core_n_1340}),
        .\reg_sbadaddr_reg[30]_2 ({core_n_1341,core_n_1342}),
        .\reg_sbadaddr_reg[30]_3 (core_n_1778),
        .\reg_sbadaddr_reg[30]_4 ({core_n_1783,core_n_1784,core_n_1785}),
        .\reg_sbadaddr_reg[30]_5 ({core_n_1788,core_n_1789}),
        .\reg_sbadaddr_reg[30]_6 ({core_n_1790,core_n_1791,core_n_1792}),
        .\reg_sbadaddr_reg[30]_7 ({core_n_1793,core_n_1794}),
        .\reg_sbadaddr_reg[30]_8 ({core_n_1795,core_n_1796}),
        .\reg_sbadaddr_reg[30]_9 ({core_n_1797,core_n_1798}),
        .\reg_sbadaddr_reg[39] (core_n_652),
        .\reg_sbadaddr_reg[39]_0 (core_n_1696),
        .\reg_sbadaddr_reg[39]_1 ({core_n_1697,core_n_1698,core_n_1699,core_n_1700}),
        .\reg_sbadaddr_reg[39]_2 ({core_n_1701,core_n_1702,core_n_1703,core_n_1704}),
        .\reg_scause_reg[0] (core_n_995),
        .\reg_scause_reg[0]_0 (core_n_1013),
        .\reg_scause_reg[1] (core_n_1010),
        .\reg_scause_reg[1]_0 (core_n_1016),
        .\reg_scause_reg[2] (wb_reg_cause),
        .\reg_scause_reg[3] (core_n_1012),
        .\reg_sepc_reg[12] (core_n_907),
        .\reg_sepc_reg[26] (core_n_1020),
        .reg_singleStepped(\csr/reg_singleStepped ),
        .\reg_sptbr_ppn_reg[0] (core_n_1001),
        .\reg_sscratch_reg[0] (core_n_977),
        .\reg_sscratch_reg[45] ({csr_io_bp_0_address[38],csr_io_bp_0_address[3:0]}),
        .\reg_sscratch_reg[45]_0 (core_n_1000),
        .\reg_sscratch_reg[59] (wb_ctrl_csr),
        .\reg_sscratch_reg[62] (_T_2518),
        .\reg_stvec_reg[32] (core_n_974),
        .\reg_stvec_reg[33] (core_n_973),
        .\reg_stvec_reg[34] (core_n_972),
        .\reg_stvec_reg[35] (core_n_971),
        .\reg_stvec_reg[36] (core_n_970),
        .\reg_stvec_reg[37] (core_n_969),
        .\reg_stvec_reg[38] (core_n_968),
        .reg_wfi_reg(core_n_1015),
        .\remainder_reg[103] ({core_n_370,core_n_371,core_n_372,core_n_373}),
        .\remainder_reg[103]_0 (core_n_375),
        .\remainder_reg[103]_1 (\remainder_reg[103] ),
        .\remainder_reg[103]_2 ({core__384_n_0,core__385_n_0,core__386_n_0,core__387_n_0}),
        .\remainder_reg[107] (\remainder_reg[107] ),
        .\remainder_reg[107]_0 (\remainder_reg[107]_0 ),
        .\remainder_reg[107]_1 ({core__380_n_0,core__381_n_0,core__382_n_0,core__383_n_0}),
        .\remainder_reg[111] (\remainder_reg[111] ),
        .\remainder_reg[111]_0 (\remainder_reg[111]_0 ),
        .\remainder_reg[111]_1 ({core__376_n_0,core__377_n_0,core__378_n_0,core__379_n_0}),
        .\remainder_reg[115] (\remainder_reg[115] ),
        .\remainder_reg[115]_0 (core_n_374),
        .\remainder_reg[115]_1 (\remainder_reg[115]_1 ),
        .\remainder_reg[115]_2 ({core__372_n_0,core__373_n_0,core__374_n_0,core__375_n_0}),
        .\remainder_reg[119] ({core_n_323,core_n_324,core_n_325,\remainder_reg[115]_0 }),
        .\remainder_reg[119]_0 ({core__368_n_0,core__369_n_0,core__370_n_0,core__371_n_0}),
        .\remainder_reg[123] ({core_n_342,core_n_343,core_n_344,core_n_345}),
        .\remainder_reg[123]_0 ({core__364_n_0,core__365_n_0,core__366_n_0,core__367_n_0}),
        .\remainder_reg[127] (core_n_327),
        .\remainder_reg[127]_0 ({core_n_328,core_n_329,core_n_330,core_n_331}),
        .\remainder_reg[127]_1 ({core_n_332,core_n_333,core_n_334,core_n_335}),
        .\remainder_reg[127]_2 ({core_n_336,core_n_337,core_n_338,core_n_339}),
        .\remainder_reg[127]_3 ({core_n_340,core_n_341}),
        .\remainder_reg[127]_4 ({core_n_346,core_n_347,core_n_348,core_n_349}),
        .\remainder_reg[127]_5 ({core_n_350,core_n_351,core_n_352,core_n_353}),
        .\remainder_reg[127]_6 (core_n_387),
        .\remainder_reg[127]_7 ({core__360_n_0,core__361_n_0,core__362_n_0,core__363_n_0}),
        .\remainder_reg[128] (core__324_n_0),
        .\remainder_reg[129] (core_n_98),
        .\remainder_reg[129]_0 (core_n_99),
        .\remainder_reg[129]_1 ({core_n_354,O,core_n_356}),
        .\remainder_reg[31] (core_n_237),
        .\remainder_reg[33] (core_n_265),
        .\remainder_reg[33]_0 (core_n_1682),
        .\remainder_reg[34] (core_n_266),
        .\remainder_reg[34]_0 (core_n_1683),
        .\remainder_reg[35] (core_n_267),
        .\remainder_reg[35]_0 (core_n_1684),
        .\remainder_reg[36] (core_n_268),
        .\remainder_reg[36]_0 (core_n_1685),
        .\remainder_reg[37] (core_n_269),
        .\remainder_reg[37]_0 (core_n_1686),
        .\remainder_reg[38] (core_n_270),
        .\remainder_reg[38]_0 (core_n_1687),
        .\remainder_reg[39] (core_n_271),
        .\remainder_reg[41] (core_n_272),
        .\remainder_reg[42] (core_n_273),
        .\remainder_reg[43] (core_n_274),
        .\remainder_reg[44] (core_n_275),
        .\remainder_reg[46] (core_n_276),
        .\remainder_reg[47] (core_n_277),
        .\remainder_reg[49] (core_n_278),
        .\remainder_reg[50] (core_n_279),
        .\remainder_reg[51] (core_n_280),
        .\remainder_reg[52] (core_n_281),
        .\remainder_reg[54] (core_n_282),
        .\remainder_reg[55] (core_n_283),
        .\remainder_reg[57] (core_n_284),
        .\remainder_reg[58] (core_n_285),
        .\remainder_reg[59] (core_n_238),
        .\remainder_reg[60] (core_n_286),
        .\remainder_reg[61] (core_n_287),
        .\remainder_reg[62] (core_n_288),
        .\remainder_reg[62]_0 ({core__664_n_0,core__665_n_0,core__666_n_0,core__667_n_0,core__668_n_0,core__669_n_0,core__670_n_0,core__671_n_0,core__672_n_0,core__673_n_0,core__674_n_0,core__675_n_0,core__676_n_0,core__677_n_0,core__678_n_0,core__679_n_0,core__680_n_0,core__681_n_0,core__682_n_0,core__683_n_0,core__684_n_0,core__685_n_0,core__686_n_0,core__687_n_0,core__688_n_0}),
        .\remainder_reg[63] (core_n_310),
        .\remainder_reg[64] ({core__351_i_2_n_0,core__351_i_3_n_0,core__351_i_4_n_0}),
        .\remainder_reg[64]_0 ({core__347_i_2_n_0,core__347_i_3_n_0,core__347_i_4_n_0,core__347_i_5_n_0}),
        .\remainder_reg[64]_1 ({core__343_i_2_n_0,core__343_i_3_n_0,core__343_i_4_n_0,core__343_i_5_n_0}),
        .\remainder_reg[64]_2 ({core__342_i_8_n_0,core__342_i_9_n_0,core__342_i_10_n_0}),
        .\remainder_reg[64]_3 (S),
        .\remainder_reg[64]_4 (\remainder_reg[64] ),
        .\remainder_reg[64]_5 (\remainder_reg[64]_0 ),
        .\remainder_reg[64]_6 ({core__357_n_0,\remainder_reg[64]_1 }),
        .\remainder_reg[64]_7 (DI),
        .\remainder_reg[64]_8 ({core__359_n_0,core__342_n_0,core__343_n_0,core__344_n_0}),
        .\remainder_reg[64]_9 (core__358_n_0),
        .\remainder_reg[65] ({core_n_105,\div/_T_103 ,core_n_107,core_n_108,core_n_109,core_n_110,core_n_111,core_n_112,core_n_113,core_n_114,core_n_115,core_n_116,core_n_117,core_n_118,core_n_119,core_n_120,core_n_121,core_n_122,core_n_123,core_n_124,core_n_125,core_n_126,core_n_127,core_n_128,core_n_129,core_n_130,core_n_131,core_n_132,core_n_133,core_n_134,core_n_135,core_n_136,core_n_137,core_n_138,core_n_139,core_n_140,core_n_141,core_n_142,core_n_143,core_n_144,core_n_145,core_n_146,core_n_147,core_n_148,core_n_149,core_n_150,core_n_151,core_n_152,core_n_153,core_n_154,core_n_155,core_n_156,core_n_157,core_n_158,core_n_159,core_n_160,core_n_161,core_n_162,core_n_163,core_n_164,core_n_165,core_n_166,core_n_167,core_n_168,core_n_169}),
        .\remainder_reg[71] ({core__416_n_0,core__417_n_0,core__418_n_0,core__419_n_0}),
        .\remainder_reg[75] ({core__412_n_0,core__413_n_0,core__414_n_0,core__415_n_0}),
        .\remainder_reg[79] ({core__408_n_0,core__409_n_0,core__410_n_0,core__411_n_0}),
        .\remainder_reg[83] ({core__404_n_0,core__405_n_0,core__406_n_0,core__407_n_0}),
        .\remainder_reg[87] ({core__400_n_0,core__401_n_0,core__402_n_0,core__403_n_0}),
        .\remainder_reg[91] ({core_n_358,core_n_359,core_n_360,core_n_361}),
        .\remainder_reg[91]_0 ({core__396_n_0,core__397_n_0,core__398_n_0,core__399_n_0}),
        .\remainder_reg[95] ({core_n_362,core_n_363,core_n_364,core_n_365}),
        .\remainder_reg[95]_0 ({core__392_n_0,core__393_n_0,core__394_n_0,core__395_n_0}),
        .\remainder_reg[99] ({core_n_366,core_n_367,core_n_368,core_n_369}),
        .\remainder_reg[99]_0 ({core__388_n_0,core__389_n_0,core__390_n_0,core__391_n_0}),
        .req_dw_reg(core_n_0),
        .\req_tag_reg[0] (dcache_n_561),
        .\req_tag_reg[0]_0 (dcache_n_562),
        .\req_tag_reg[1] (dcache_n_563),
        .\req_tag_reg[1]_0 (dcache_n_565),
        .\req_tag_reg[1]_1 (dcache_n_560),
        .\req_tag_reg[1]_2 (dcache_n_564),
        .\req_tag_reg[1]_3 (dcache_n_566),
        .\req_tag_reg[1]_4 (dcache_n_559),
        .\req_tag_reg[4] (frontend_n_416),
        .resHi_reg(core_n_104),
        .resp_valid_0_reg(ptw_n_184),
        .resp_valid_1_reg(s2_valid_reg),
        .\s1_pc_reg[1] (core_n_1029),
        .\s1_pc_reg[26] (frontend_n_126),
        .\s1_pc_reg[31] (frontend_n_152),
        .\s1_pc_reg[39] (core_n_651),
        .\s1_pc_reg[39]_0 (frontend_io_cpu_req_bits_pc),
        .\s1_pc_reg[39]_1 ({core_n_1430,core_n_1431,core_n_1432,core_n_1433}),
        .\s1_pc_reg[39]_2 ({core_n_1434,core_n_1435,core_n_1436,core_n_1437}),
        .\s1_pc_reg[39]_3 ({core_n_1438,core_n_1439,core_n_1440,core_n_1441}),
        .\s1_pc_reg[39]_4 ({core_n_1442,core_n_1443,core_n_1444,core_n_1445}),
        .\s1_pc_reg[39]_5 (core_n_1705),
        .\s1_pc_reg[39]_6 ({s1_pc[39:38],s1_pc[11:2]}),
        .\s1_pc_reg[4] (\csr/reg_stvec ),
        .\s1_pc_reg[4]_0 (\csr/reg_mtvec ),
        .\s1_pc_reg[5] (core_n_1011),
        .\s1_req_addr_reg[2] (ptw_n_137),
        .\s1_req_addr_reg[2]_0 (ptw_n_152),
        .\s1_req_addr_reg[2]_1 (ptw_n_148),
        .\s1_req_addr_reg[2]_2 (ptw_n_155),
        .\s1_req_addr_reg[31] ({dcache_n_140,dcache_n_141,dcache_n_145,dcache_n_147,dcache_n_151,dcache_n_153,dcache_n_159,_T_1701[2:0],_T_628}),
        .\s1_req_addr_reg[39] ({_T_2770[24:21],_T_2770[19:18],_T_2770[16:15],_T_2770[13:10],_T_2770[8:7],_T_2770[5:2],_T_2770[0]}),
        .\s1_req_addr_reg[39]_0 ({core_n_1608,core_n_1609,core_n_1610,core_n_1611}),
        .\s1_req_addr_reg[39]_1 ({core_n_1612,core_n_1613,core_n_1614,core_n_1615}),
        .\s1_req_addr_reg[39]_2 ({core_n_1688,core_n_1689,core_n_1690,core_n_1691}),
        .\s1_req_addr_reg[39]_3 ({core_n_1692,core_n_1693,core_n_1694,core_n_1695}),
        .\s1_req_addr_reg[39]_4 (core_n_1787),
        .\s1_req_addr_reg[3] (core_n_1786),
        .\s1_req_cmd_reg[4] (dcacheArb_io_requestor_1_req_bits_cmd),
        .s1_req_phys_reg(dcache_n_89),
        .s1_req_phys_reg_0(dcache_n_584),
        .\s1_req_typ_reg[0] (dcache_n_615),
        .\s1_req_typ_reg[0]_0 (dcache_n_429),
        .\s1_req_typ_reg[0]_1 (dcache_n_617),
        .\s1_req_typ_reg[0]_2 (dcache_n_624),
        .\s1_req_typ_reg[0]_3 (dcache_n_619),
        .\s1_req_typ_reg[1] (dcache_n_621),
        .s1_valid_reg(core_n_647),
        .\s2_pc_reg[1] (s2_pc[1]),
        .s2_replay(s2_replay),
        .\s2_req_addr_reg[31] (dcache_io_ptw_status_dprv),
        .\s2_req_cmd_reg[1] (dcache_n_369),
        .\s2_req_tag_reg[5] (dcache_n_541),
        .\s2_req_tag_reg[5]_0 (dcache_n_554),
        .\s2_req_tag_reg[6] (dcacheArb_io_requestor_1_resp_bits_tag),
        .\s2_req_tag_reg[6]_0 (dcache_n_552),
        .\s2_req_typ_reg[0] (_GEN_274[29:10]),
        .s2_tlb_resp_cacheable_reg(core_n_752),
        .s2_valid_reg(core_n_749),
        .shamt(\alu/shamt ),
        .\state_reg[0] (core__192_n_0),
        .\state_reg[0]_0 (ptw_n_2),
        .\state_reg[0]_1 (ptw_n_52),
        .\state_reg[0]_2 (core__184_n_0),
        .\state_reg[1] (core_n_1028),
        .\state_reg[1]_0 (core__191_n_0),
        .\state_reg[1]_1 (ptw_n_1),
        .\state_reg[2] (core_n_101),
        .sys_reset_reg(core__501_n_0),
        .sys_reset_reg_0(core__716_n_0),
        .sys_reset_reg_1(core__503_n_0),
        .sys_reset_reg_2(core__502_n_0),
        .target_reset(target_reset),
        .tile_auto_int_sync_xing_sinklzy_in_0_sync_0(tile_auto_int_sync_xing_sinklzy_in_0_sync_0),
        .tile_auto_int_sync_xing_sinklzy_in_0_sync_1(tile_auto_int_sync_xing_sinklzy_in_0_sync_1),
        .tile_auto_int_sync_xing_sinklzy_in_1_sync_0(tile_auto_int_sync_xing_sinklzy_in_1_sync_0),
        .tile_auto_int_sync_xing_sinklzy_in_2_sync_0(tile_auto_int_sync_xing_sinklzy_in_2_sync_0),
        .tlb_io_req_bits_sfence_bits_rs2(tlb_io_req_bits_sfence_bits_rs2),
        .\trig_jalr_count_reg[0]_0 (core_n_1365),
        .\trig_jalr_count_reg[0]_1 ({core_n_1469,core_n_1470,core_n_1471,core_n_1472}),
        .\trig_jalr_count_reg[0]_2 ({core_n_1473,core_n_1474,core_n_1475,core_n_1476}),
        .\trig_jalr_count_reg[0]_3 ({core_n_1477,core_n_1478,core_n_1479,core_n_1480}),
        .\trig_jalr_count_reg[0]_4 ({core_n_1481,core_n_1482,core_n_1483,core_n_1484}),
        .\trig_jalr_count_reg[0]_5 ({core_n_1485,core_n_1486,core_n_1487,core_n_1488}),
        .\trig_jalr_count_reg[0]_6 (core_n_1489),
        .\trig_mem_data_reg[126]_0 ({_GEN_277[126],_GEN_277[62]}),
        .\trig_mem_data_reg[127]_0 (trigB),
        .\trig_mem_data_reg[63]_0 (trigA),
        .\trig_pc_reg[0]_0 (core_n_30),
        .\trig_pc_reg[0]_1 (core_n_1349),
        .\trig_pc_reg[0]_2 ({core_n_1490,core_n_1491,core_n_1492,core_n_1493}),
        .\trig_pc_reg[0]_3 ({core_n_1591,core_n_1592,core_n_1593,core_n_1594}),
        .\trig_pc_reg[0]_4 ({core_n_1595,core_n_1596,core_n_1597,core_n_1598}),
        .\trig_pc_reg[0]_5 ({core_n_1599,core_n_1600,core_n_1601,core_n_1602}),
        .\trig_pc_reg[0]_6 ({core_n_1603,core_n_1604,core_n_1605,core_n_1606}),
        .\trig_pc_reg[0]_7 (core_n_1607),
        .\trig_pc_reg[63]_0 ({core_n_1494,core_n_1495,core_n_1496,core_n_1497,core_n_1498,core_n_1499,core_n_1500,core_n_1501,core_n_1502,core_n_1503,core_n_1504,core_n_1505,core_n_1506,core_n_1507,core_n_1508,core_n_1509,core_n_1510,core_n_1511,core_n_1512,core_n_1513,core_n_1514,core_n_1515,core_n_1516,core_n_1517,core_n_1518,core_n_1519,core_n_1520,core_n_1521,core_n_1522,core_n_1523,core_n_1524,core_n_1525,core_n_1526,core_n_1527,core_n_1528,core_n_1529,core_n_1530,core_n_1531,core_n_1532,core_n_1533,core_n_1534,core_n_1535,core_n_1536,core_n_1537,core_n_1538,core_n_1539,core_n_1540,core_n_1541,core_n_1542,core_n_1543,core_n_1544,core_n_1545,core_n_1546,core_n_1547,core_n_1548,core_n_1549,core_n_1550,core_n_1551,core_n_1552,core_n_1553,core_n_1554,core_n_1555,core_n_1556,core_n_1557}),
        .\trig_pc_reg[63]_1 (_T_1944),
        .trig_pc_valid_reg_0(core_n_1350),
        .trig_pc_valid_reg_1(core__434_n_0),
        .trig_pc_valid_reg_2(core__266_n_0),
        .\trig_state_reg[0]_0 (core_n_1346),
        .\trig_state_reg[0]_1 (core__265_n_0),
        .\trig_state_reg[1]_0 (core_n_1345),
        .\trig_state_reg[1]_1 (core_n_1347),
        .\trig_state_reg[1]_2 (core_n_1348),
        .\trig_state_reg[1]_3 ({core_n_1446,core_n_1447,core_n_1448,core_n_1449}),
        .\trig_state_reg[1]_4 ({core_n_1452,core_n_1453,core_n_1454,core_n_1455}),
        .\trig_state_reg[1]_5 ({core_n_1456,core_n_1457,core_n_1458,core_n_1459}),
        .\trig_state_reg[1]_6 ({core_n_1460,core_n_1461,core_n_1462,core_n_1463}),
        .\trig_state_reg[1]_7 ({core_n_1464,core_n_1465,core_n_1466,core_n_1467}),
        .\trig_state_reg[1]_8 (core_n_1468),
        .\valid_reg[0] (core_n_1839),
        .\valid_reg[0]_0 (dcache_n_634),
        .\valid_reg[1] (core_n_686),
        .\valid_reg[1]_0 (dcache_n_633),
        .\valid_reg[2] (dcache_n_134),
        .\valid_reg[3] (core_n_551),
        .\valid_reg[3]_0 (core_n_682),
        .\valid_reg[3]_1 (frontend_io_cpu_sfence_bits_rs1),
        .\valid_reg[3]_2 (\tlb/_GEN_29 ),
        .\valid_reg[3]_3 (core_n_685),
        .\valid_reg[3]_4 (\tlb/_T_815 ),
        .\valid_reg[4] (dcache_n_133),
        .\wb_ctrl_csr_reg[0]_0 (core__121_n_0),
        .\wb_ctrl_csr_reg[0]_1 (core__510_n_0),
        .\wb_ctrl_csr_reg[0]_10 (core__550_n_0),
        .\wb_ctrl_csr_reg[0]_2 (core__460_n_0),
        .\wb_ctrl_csr_reg[0]_3 (\csr/p_1_in ),
        .\wb_ctrl_csr_reg[0]_4 (core__504_n_0),
        .\wb_ctrl_csr_reg[0]_5 ({core__505_n_0,core__506_n_0,core__507_n_0,core__508_n_0,core__509_n_0}),
        .\wb_ctrl_csr_reg[0]_6 (core__598_n_0),
        .\wb_ctrl_csr_reg[0]_7 (core__551_n_0),
        .\wb_ctrl_csr_reg[0]_8 ({core__552_n_0,core__553_n_0,core__554_n_0,core__555_n_0,core__556_n_0,core__557_n_0}),
        .\wb_ctrl_csr_reg[0]_9 (core__558_n_0),
        .\wb_ctrl_csr_reg[2]_0 (core__125_n_0),
        .wb_ctrl_div(wb_ctrl_div),
        .wb_ctrl_fence_i_reg_0(core_n_28),
        .wb_ctrl_mem(wb_ctrl_mem),
        .wb_ctrl_mem_reg_0(dcache_n_557),
        .wb_ctrl_wxd(wb_ctrl_wxd),
        .\wb_reg_cause_reg[0]_0 (core_n_1320),
        .\wb_reg_cause_reg[0]_1 ({core_n_2151,core_n_2152,core_n_2153,core_n_2154}),
        .\wb_reg_cause_reg[0]_10 ({core_n_2184,core_n_2185,core_n_2186,core_n_2187}),
        .\wb_reg_cause_reg[0]_11 ({core_n_2188,core_n_2189,core_n_2190,core_n_2191}),
        .\wb_reg_cause_reg[0]_12 ({core_n_2192,core_n_2193,core_n_2194,core_n_2195}),
        .\wb_reg_cause_reg[0]_13 ({core_n_2196,core_n_2197,core_n_2198}),
        .\wb_reg_cause_reg[0]_14 ({core_n_2199,core_n_2200,core_n_2201}),
        .\wb_reg_cause_reg[0]_2 ({core_n_2155,core_n_2156,core_n_2157,core_n_2158}),
        .\wb_reg_cause_reg[0]_3 ({core_n_2159,core_n_2160,core_n_2161,core_n_2162}),
        .\wb_reg_cause_reg[0]_4 (core_n_2163),
        .\wb_reg_cause_reg[0]_5 ({core_n_2164,core_n_2165,core_n_2166,core_n_2167}),
        .\wb_reg_cause_reg[0]_6 ({core_n_2168,core_n_2169,core_n_2170,core_n_2171}),
        .\wb_reg_cause_reg[0]_7 ({core_n_2172,core_n_2173,core_n_2174,core_n_2175}),
        .\wb_reg_cause_reg[0]_8 ({core_n_2176,core_n_2177,core_n_2178,core_n_2179}),
        .\wb_reg_cause_reg[0]_9 ({core_n_2180,core_n_2181,core_n_2182,core_n_2183}),
        .\wb_reg_cause_reg[2]_0 (core__433_n_0),
        .\wb_reg_cause_reg[3]_0 (mem_reg_cause),
        .\wb_reg_cause_reg[63]_0 (dcache_n_558),
        .\wb_reg_cause_reg[63]_1 (_T_2499),
        .\wb_reg_cause_reg[63]_2 (_T_2434),
        .\wb_reg_cause_reg[63]_3 (_T_2425),
        .\wb_reg_cause_reg[63]_4 (_T_2431),
        .\wb_reg_cause_reg[63]_5 (_T_2428),
        .\wb_reg_cause_reg[63]_6 (_T_2498),
        .\wb_reg_inst_reg[21]_0 (core__108_n_0),
        .\wb_reg_inst_reg[21]_1 (core__106_n_0),
        .\wb_reg_inst_reg[21]_2 (core__113_n_0),
        .\wb_reg_inst_reg[21]_3 (core__110_n_0),
        .\wb_reg_inst_reg[21]_4 (core__109_n_0),
        .\wb_reg_inst_reg[21]_5 (core__122_n_0),
        .\wb_reg_inst_reg[22]_0 (core__105_n_0),
        .\wb_reg_inst_reg[22]_1 (core__119_n_0),
        .\wb_reg_inst_reg[26]_0 (core__123_n_0),
        .\wb_reg_inst_reg[29]_0 (core__112_n_0),
        .\wb_reg_inst_reg[29]_1 (core__114_n_0),
        .\wb_reg_inst_reg[30]_0 (core__124_n_0),
        .\wb_reg_inst_reg[30]_1 (core__115_n_0),
        .\wb_reg_inst_reg[31]_0 ({_T_20810,core_n_1104,core_n_1105,core_n_1106,core_n_1107,core_n_1108,core_n_1109,core_n_1110,core_n_1111,core_n_1112,core_n_1113,core_n_1114,core_n_1115,core_n_1116,core_n_1117,core_n_1118,core_n_1119,core_n_1120,core_n_1121,core_n_1122,mem_waddr}),
        .\wb_reg_inst_reg[7]_0 (frontend_n_365),
        .\wb_reg_inst_reg[7]_1 (frontend_n_351),
        .\wb_reg_inst_reg[9]_0 (core__318_n_0),
        .\wb_reg_inst_reg[9]_1 (core__317_n_0),
        .\wb_reg_inst_reg[9]_2 (core__316_n_0),
        .\wb_reg_inst_reg[9]_3 (core__319_n_0),
        .\wb_reg_pc_reg[34]_0 ({mem_reg_pc[34:32],core_n_1354}),
        .\wb_reg_pc_reg[39]_0 ({mem_reg_pc[39:35],mem_reg_pc[31],mem_reg_pc[27:1]}),
        .\wb_reg_pc_reg[39]_1 (\csr/_GEN_350 ),
        .\wb_reg_pc_reg[39]_2 (\csr/_GEN_364 ),
        .\wb_reg_pc_reg[39]_3 (\csr/_GEN_369 ),
        .wb_reg_replay(wb_reg_replay),
        .wb_reg_replay_reg_0(dcache_n_555),
        .wb_reg_replay_reg_1(dcache_n_556),
        .wb_reg_replay_reg_2(core__186_n_0),
        .wb_reg_valid(wb_reg_valid),
        .wb_reg_valid_reg_0(core__118_n_0),
        .wb_reg_xcpt(wb_reg_xcpt));
  LUT4 #(
    .INIT(16'hE200)) 
    core__10
       (.I0(_GEN_274[60]),
        .I1(frontend_n_351),
        .I2(_T_1406[60]),
        .I3(frontend_n_352),
        .O(core__10_n_0));
  LUT4 #(
    .INIT(16'h00E2)) 
    core__100
       (.I0(frontend_io_cpu_resp_bits_pc[1]),
        .I1(\ibuf/_T_100 ),
        .I2(core_n_1088),
        .I3(csr_io_bp_0_address[1]),
        .O(core__100_n_0));
  LUT5 #(
    .INIT(32'h0000B847)) 
    core__101
       (.I0(core_n_1088),
        .I1(\ibuf/_T_100 ),
        .I2(frontend_io_cpu_resp_bits_pc[1]),
        .I3(csr_io_bp_0_address[1]),
        .I4(csr_io_bp_0_address[0]),
        .O(core__101_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2487" *) 
  LUT5 #(
    .INIT(32'h40444444)) 
    core__102
       (.I0(csr_io_status_debug),
        .I1(\csr/reg_dcsr_step ),
        .I2(\csr/reg_singleStepped ),
        .I3(dcache_n_555),
        .I4(core_n_1015),
        .O(core__102_n_0));
  LUT4 #(
    .INIT(16'h5C55)) 
    core__103
       (.I0(core_n_82),
        .I1(\csr/_T_4899 [6]),
        .I2(core_n_894),
        .I3(core_n_895),
        .O(core__103_n_0));
  LUT4 #(
    .INIT(16'h5C55)) 
    core__104
       (.I0(\csr/_T_286__0 ),
        .I1(\csr/_T_4899 [6]),
        .I2(core__108_n_0),
        .I3(core_n_896),
        .O(core__104_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2489" *) 
  LUT4 #(
    .INIT(16'hDFFF)) 
    core__105
       (.I0(csr_io_rw_addr[2]),
        .I1(core__124_n_0),
        .I2(csr_io_rw_addr[0]),
        .I3(csr_io_rw_addr[1]),
        .O(core__105_n_0));
  LUT5 #(
    .INIT(32'hFFF7FFFF)) 
    core__106
       (.I0(csr_io_rw_addr[1]),
        .I1(csr_io_rw_addr[0]),
        .I2(csr_io_rw_addr[2]),
        .I3(core_n_977),
        .I4(core_n_957),
        .O(core__106_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    core__107
       (.I0(\csr/_T_5074 ),
        .I1(csr_io_status_debug),
        .O(core__107_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2561" *) 
  LUT2 #(
    .INIT(4'hB)) 
    core__108
       (.I0(core_n_997),
        .I1(csr_io_rw_addr[1]),
        .O(core__108_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2561" *) 
  LUT2 #(
    .INIT(4'hB)) 
    core__109
       (.I0(core_n_1000),
        .I1(csr_io_rw_addr[1]),
        .O(core__109_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__11
       (.I0(_GEN_274[59]),
        .I1(frontend_n_351),
        .I2(_T_1406[59]),
        .I3(frontend_n_352),
        .O(core__11_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2489" *) 
  LUT4 #(
    .INIT(16'hEFFF)) 
    core__110
       (.I0(core__112_n_0),
        .I1(csr_io_rw_addr[1]),
        .I2(csr_io_rw_addr[0]),
        .I3(csr_io_rw_addr[2]),
        .O(core__110_n_0));
  LUT5 #(
    .INIT(32'h22F2FFFF)) 
    core__111
       (.I0(frontend_io_ptw_pmp_5_addr[20]),
        .I1(core__122_n_0),
        .I2(frontend_io_ptw_pmp_2_addr[20]),
        .I3(core_n_996),
        .I4(core_n_994),
        .O(core__111_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    core__112
       (.I0(csr_io_rw_addr[9]),
        .I1(csr_io_rw_addr[10]),
        .I2(csr_io_rw_addr[7]),
        .I3(core_n_999),
        .I4(csr_io_rw_addr[11]),
        .I5(core_n_1001),
        .O(core__112_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2498" *) 
  LUT4 #(
    .INIT(16'hEFFF)) 
    core__113
       (.I0(core__114_n_0),
        .I1(csr_io_rw_addr[1]),
        .I2(csr_io_rw_addr[0]),
        .I3(csr_io_rw_addr[2]),
        .O(core__113_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    core__114
       (.I0(csr_io_rw_addr[9]),
        .I1(csr_io_rw_addr[10]),
        .I2(csr_io_rw_addr[7]),
        .I3(core_n_999),
        .I4(csr_io_rw_addr[11]),
        .I5(core_n_1001),
        .O(core__114_n_0));
  LUT3 #(
    .INIT(8'h20)) 
    core__115
       (.I0(core_n_1003),
        .I1(csr_io_rw_addr[10]),
        .I2(csr_io_rw_addr[9]),
        .O(core__115_n_0));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    core__116
       (.I0(\csr/reg_mtvec ),
        .I1(core_n_1004),
        .I2(\csr/reg_stvec ),
        .I3(core_n_1011),
        .I4(core__433_n_0),
        .I5(core_n_1009),
        .O(core__116_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2556" *) 
  LUT3 #(
    .INIT(8'h04)) 
    core__117
       (.I0(core_n_1004),
        .I1(core_n_1009),
        .I2(core_n_1015),
        .O(core__117_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2556" *) 
  LUT2 #(
    .INIT(4'hB)) 
    core__118
       (.I0(core_n_1003),
        .I1(core_n_1009),
        .O(core__118_n_0));
  LUT6 #(
    .INIT(64'hAAAAAA88AAAAAA8B)) 
    core__119
       (.I0(core_n_1013),
        .I1(csr_io_rw_addr[2]),
        .I2(csr_io_rw_addr[0]),
        .I3(csr_io_rw_addr[1]),
        .I4(core__121_n_0),
        .I5(frontend_io_ptw_status_prv[0]),
        .O(core__119_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__12
       (.I0(_GEN_274[58]),
        .I1(frontend_n_351),
        .I2(_T_1406[58]),
        .I3(frontend_n_352),
        .O(core__12_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2487" *) 
  LUT2 #(
    .INIT(4'h1)) 
    core__120
       (.I0(csr_io_status_debug),
        .I1(core_n_1015),
        .O(core__120_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2497" *) 
  LUT4 #(
    .INIT(16'hEFFF)) 
    core__121
       (.I0(wb_ctrl_csr[0]),
        .I1(wb_ctrl_csr[1]),
        .I2(wb_ctrl_csr[2]),
        .I3(wb_reg_valid),
        .O(core__121_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2498" *) 
  LUT4 #(
    .INIT(16'hEFFF)) 
    core__122
       (.I0(core__124_n_0),
        .I1(csr_io_rw_addr[1]),
        .I2(csr_io_rw_addr[0]),
        .I3(csr_io_rw_addr[2]),
        .O(core__122_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2490" *) 
  LUT4 #(
    .INIT(16'hFBFF)) 
    core__123
       (.I0(csr_io_rw_addr[6]),
        .I1(csr_io_rw_addr[10]),
        .I2(core_n_1018),
        .I3(csr_io_rw_addr[4]),
        .O(core__123_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2490" *) 
  LUT4 #(
    .INIT(16'hFEFF)) 
    core__124
       (.I0(csr_io_rw_addr[10]),
        .I1(csr_io_rw_addr[6]),
        .I2(core_n_1018),
        .I3(csr_io_rw_addr[4]),
        .O(core__124_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2497" *) 
  LUT4 #(
    .INIT(16'h4000)) 
    core__125
       (.I0(wb_ctrl_csr[2]),
        .I1(wb_reg_valid),
        .I2(wb_ctrl_csr[0]),
        .I3(wb_ctrl_csr[1]),
        .O(core__125_n_0));
  LUT3 #(
    .INIT(8'h45)) 
    core__126
       (.I0(frontend_io_ptw_status_prv[1]),
        .I1(core_n_85),
        .I2(frontend_io_ptw_status_prv[0]),
        .O(core__126_n_0));
  LUT6 #(
    .INIT(64'hF999999999999999)) 
    core__127
       (.I0(csr_io_bp_0_address[3]),
        .I1(core_n_1330),
        .I2(csr_io_bp_0_address[1]),
        .I3(csr_io_bp_0_control_tmatch),
        .I4(csr_io_bp_0_address[0]),
        .I5(csr_io_bp_0_address[2]),
        .O(core__127_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    core__128
       (.I0(\bpu/_T_134 ),
        .I1(csr_io_bp_0_control_action),
        .O(core__128_n_0));
  CARRY4 core__128_i_14
       (.CI(core__128_i_28_n_0),
        .CO({core__128_i_14_n_0,core__128_i_14_n_1,core__128_i_14_n_2,core__128_i_14_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_2121,core_n_2122,core_n_2123,core_n_2124}));
  CARRY4 core__128_i_19
       (.CI(core__128_i_33_n_0),
        .CO({core__128_i_19_n_0,core__128_i_19_n_1,core__128_i_19_n_2,core__128_i_19_n_3}),
        .CYINIT(\<const0> ),
        .DI({core_n_2125,core_n_2126,core_n_2127,core_n_2128}),
        .S({core_n_2129,core_n_2130,core_n_2131,core_n_2132}));
  CARRY4 core__128_i_2
       (.CI(core__128_i_4_n_0),
        .CO(\bpu/_T_132 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,core_n_2102}));
  CARRY4 core__128_i_28
       (.CI(\<const0> ),
        .CO({core__128_i_28_n_0,core__128_i_28_n_1,core__128_i_28_n_2,core__128_i_28_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_2141,core_n_2142,core_n_2143,core_n_2144}));
  CARRY4 core__128_i_3
       (.CI(core__128_i_6_n_0),
        .CO({\bpu/_T_105 ,core__128_i_3_n_1,core__128_i_3_n_2,core__128_i_3_n_3}),
        .CYINIT(\<const0> ),
        .DI({core__717_n_0,core_n_2103,core_n_2104,core_n_2105}),
        .S({frontend_n_92,core_n_2106,core_n_2107,core_n_2108}));
  CARRY4 core__128_i_33
       (.CI(core__128_i_46_n_0),
        .CO({core__128_i_33_n_0,core__128_i_33_n_1,core__128_i_33_n_2,core__128_i_33_n_3}),
        .CYINIT(\<const0> ),
        .DI({core_n_2133,core_n_2134,core_n_2135,core_n_2136}),
        .S({core_n_2137,core_n_2138,core_n_2139,core_n_2140}));
  CARRY4 core__128_i_4
       (.CI(core__128_i_14_n_0),
        .CO({core__128_i_4_n_0,core__128_i_4_n_1,core__128_i_4_n_2,core__128_i_4_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_2109,core_n_2110,core_n_2111,core_n_2112}));
  CARRY4 core__128_i_46
       (.CI(\<const0> ),
        .CO({core__128_i_46_n_0,core__128_i_46_n_1,core__128_i_46_n_2,core__128_i_46_n_3}),
        .CYINIT(\<const1> ),
        .DI({core_n_2145,core_n_2146,core_n_2147,core__100_n_0}),
        .S({core_n_2148,core_n_2149,core_n_2150,core__101_n_0}));
  CARRY4 core__128_i_6
       (.CI(core__128_i_19_n_0),
        .CO({core__128_i_6_n_0,core__128_i_6_n_1,core__128_i_6_n_2,core__128_i_6_n_3}),
        .CYINIT(\<const0> ),
        .DI({core_n_2113,core_n_2114,core_n_2115,core_n_2116}),
        .S({core_n_2117,core_n_2118,core_n_2119,core_n_2120}));
  LUT6 #(
    .INIT(64'h00000000F4A45404)) 
    core__129
       (.I0(frontend_io_ptw_status_prv[1]),
        .I1(csr_io_bp_0_control_u),
        .I2(frontend_io_ptw_status_prv[0]),
        .I3(csr_io_bp_0_control_s),
        .I4(csr_io_bp_0_control_m),
        .I5(csr_io_status_debug),
        .O(core__129_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__13
       (.I0(_GEN_274[57]),
        .I1(frontend_n_351),
        .I2(_T_1406[57]),
        .I3(frontend_n_352),
        .O(core__13_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__130
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2284),
        .I3(core_n_2204),
        .I4(dcacheArb_io_requestor_1_req_bits_addr[33]),
        .O(core__130_n_0));
  CARRY4 core__130_i_4
       (.CI(core__161_i_1_n_0),
        .CO({core__130_i_4_n_0,core__130_i_4_n_1,core__130_i_4_n_2,core__130_i_4_n_3}),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[35:32]),
        .O(dcacheArb_io_requestor_1_req_bits_addr[35:32]),
        .S({core__288_n_0,core__287_n_0,core_rep__13_n_0,core__286_n_0}));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__131
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2282),
        .I3(core_n_2205),
        .I4(dcacheArb_io_requestor_1_req_bits_addr[34]),
        .O(core__131_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__132
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2280),
        .I3(core_n_2206),
        .I4(dcacheArb_io_requestor_1_req_bits_addr[35]),
        .O(core__132_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__133
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2279),
        .I3(core_n_2207),
        .I4(dcacheArb_io_requestor_1_req_bits_addr[36]),
        .O(core__133_n_0));
  CARRY4 core__133_i_3
       (.CI(core__130_i_4_n_0),
        .CO({core__133_i_3_n_0,core__133_i_3_n_1,core__133_i_3_n_2,core__133_i_3_n_3}),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[39:36]),
        .O({alu_io_adder_out,dcacheArb_io_requestor_1_req_bits_addr[38:36]}),
        .S({core_rep__15_n_0,core__290_n_0,core__289_n_0,core_rep__14_n_0}));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__134
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2277),
        .I3(core_n_2208),
        .I4(dcacheArb_io_requestor_1_req_bits_addr[37]),
        .O(core__134_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__135
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2275),
        .I3(core_n_2209),
        .I4(dcacheArb_io_requestor_1_req_bits_addr[38]),
        .O(core__135_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__136
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2273),
        .I3(core_n_2210),
        .I4(alu_io_adder_out),
        .O(core__136_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__137
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2271),
        .I3(core_n_2211),
        .I4(core__137_i_3_n_7),
        .O(core__137_n_0));
  CARRY4 core__137_i_3
       (.CI(core__133_i_3_n_0),
        .CO({core__137_i_3_n_0,core__137_i_3_n_1,core__137_i_3_n_2,core__137_i_3_n_3}),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[43:40]),
        .O({core__137_i_3_n_4,core__137_i_3_n_5,core__137_i_3_n_6,core__137_i_3_n_7}),
        .S({core__305_n_0,core_rep__16_n_0,core__267_n_0,core__307_n_0}));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__138
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2269),
        .I3(core_n_2212),
        .I4(core__137_i_3_n_6),
        .O(core__138_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__139
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2267),
        .I3(core_n_2213),
        .I4(core__137_i_3_n_5),
        .O(core__139_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__14
       (.I0(_GEN_274[56]),
        .I1(frontend_n_351),
        .I2(_T_1406[56]),
        .I3(frontend_n_352),
        .O(core__14_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__140
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2265),
        .I3(core_n_2214),
        .I4(core__137_i_3_n_4),
        .O(core__140_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__141
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2263),
        .I3(core_n_2215),
        .I4(core__141_i_3_n_7),
        .O(core__141_n_0));
  CARRY4 core__141_i_3
       (.CI(core__137_i_3_n_0),
        .CO({core__141_i_3_n_0,core__141_i_3_n_1,core__141_i_3_n_2,core__141_i_3_n_3}),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[47:44]),
        .O({core__141_i_3_n_4,core__141_i_3_n_5,core__141_i_3_n_6,core__141_i_3_n_7}),
        .S({core__304_n_0,core__303_n_0,core_rep__17_n_0,core__306_n_0}));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__142
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2261),
        .I3(core_n_2216),
        .I4(core__141_i_3_n_6),
        .O(core__142_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__143
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2259),
        .I3(core_n_2217),
        .I4(core__141_i_3_n_5),
        .O(core__143_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__144
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2256),
        .I3(core_n_2218),
        .I4(core__141_i_3_n_4),
        .O(core__144_n_0));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__145
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2254),
        .I3(core_n_2318),
        .I4(core_n_2223),
        .I5(core__145_i_4_n_7),
        .O(core__145_n_0));
  CARRY4 core__145_i_4
       (.CI(core__141_i_3_n_0),
        .CO({core__145_i_4_n_0,core__145_i_4_n_1,core__145_i_4_n_2,core__145_i_4_n_3}),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[51:48]),
        .O({core__145_i_4_n_4,core__145_i_4_n_5,core__145_i_4_n_6,core__145_i_4_n_7}),
        .S({core_rep__19_n_0,core__302_n_0,core__301_n_0,core_rep__18_n_0}));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__146
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2253),
        .I3(core_n_2319),
        .I4(core_n_2224),
        .I5(core__145_i_4_n_6),
        .O(core__146_n_0));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__147
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2252),
        .I3(core_n_2320),
        .I4(core_n_2225),
        .I5(core__145_i_4_n_5),
        .O(core__147_n_0));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__148
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2251),
        .I3(core_n_2321),
        .I4(core_n_2226),
        .I5(core__145_i_4_n_4),
        .O(core__148_n_0));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__149
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2250),
        .I3(core_n_2322),
        .I4(core_n_2227),
        .I5(core__149_i_4_n_7),
        .O(core__149_n_0));
  CARRY4 core__149_i_4
       (.CI(core__145_i_4_n_0),
        .CO({core__149_i_4_n_0,core__149_i_4_n_1,core__149_i_4_n_2,core__149_i_4_n_3}),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[55:52]),
        .O({core__149_i_4_n_4,core__149_i_4_n_5,core__149_i_4_n_6,core__149_i_4_n_7}),
        .S({core__297_n_0,core_rep__20_n_0,core__300_n_0,core__299_n_0}));
  LUT4 #(
    .INIT(16'hE200)) 
    core__15
       (.I0(_GEN_274[55]),
        .I1(frontend_n_351),
        .I2(_T_1406[55]),
        .I3(frontend_n_352),
        .O(core__15_n_0));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__150
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2249),
        .I3(core_n_2323),
        .I4(core_n_2228),
        .I5(core__149_i_4_n_6),
        .O(core__150_n_0));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__151
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2248),
        .I3(core_n_2324),
        .I4(core_n_2229),
        .I5(core__149_i_4_n_5),
        .O(core__151_n_0));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__152
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2247),
        .I3(core_n_2325),
        .I4(core_n_2230),
        .I5(core__149_i_4_n_4),
        .O(core__152_n_0));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__153
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2246),
        .I3(core_n_2326),
        .I4(core_n_2231),
        .I5(core__153_i_4_n_7),
        .O(core__153_n_0));
  CARRY4 core__153_i_4
       (.CI(core__149_i_4_n_0),
        .CO({core__153_i_4_n_0,core__153_i_4_n_1,core__153_i_4_n_2,core__153_i_4_n_3}),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[59:56]),
        .O({core__153_i_4_n_4,core__153_i_4_n_5,core__153_i_4_n_6,core__153_i_4_n_7}),
        .S({core__296_n_0,core__295_n_0,core_rep__21_n_0,core__298_n_0}));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__154
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2245),
        .I3(core_n_2327),
        .I4(core_n_2232),
        .I5(core__153_i_4_n_6),
        .O(core__154_n_0));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__155
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2244),
        .I3(core_n_2328),
        .I4(core_n_2233),
        .I5(core__153_i_4_n_5),
        .O(core__155_n_0));
  LUT6 #(
    .INIT(64'hAAAA8AAA22220222)) 
    core__156
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2243),
        .I3(core_n_2329),
        .I4(core_n_2234),
        .I5(core__153_i_4_n_4),
        .O(core__156_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__157
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2242),
        .I3(core_n_2219),
        .I4(core__157_i_3_n_7),
        .O(core__157_n_0));
  CARRY4 core__157_i_3
       (.CI(core__153_i_4_n_0),
        .CO({core__157_i_3_n_1,core__157_i_3_n_2,core__157_i_3_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,alu_io_in1[62:60]}),
        .O({core__157_i_3_n_4,core__157_i_3_n_5,core__157_i_3_n_6,core__157_i_3_n_7}),
        .S({core__292_n_0,core__294_n_0,core__293_n_0,core_rep__22_n_0}));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__158
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2241),
        .I3(core_n_2220),
        .I4(core__157_i_3_n_6),
        .O(core__158_n_0));
  LUT5 #(
    .INIT(32'h8AAA0222)) 
    core__159
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2240),
        .I3(core_n_2221),
        .I4(core__157_i_3_n_5),
        .O(core__159_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__16
       (.I0(_GEN_274[54]),
        .I1(frontend_n_351),
        .I2(_T_1406[54]),
        .I3(frontend_n_352),
        .O(core__16_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2496" *) 
  LUT4 #(
    .INIT(16'hA820)) 
    core__160
       (.I0(core_n_0),
        .I1(\alu/_T_217 ),
        .I2(core_n_2222),
        .I3(core__157_i_3_n_4),
        .O(core__160_n_0));
  LUT5 #(
    .INIT(32'h000088A0)) 
    core__161
       (.I0(mem_ctrl_fp),
        .I1(dcacheArb_io_requestor_1_req_bits_addr[31]),
        .I2(core_n_2203),
        .I3(\alu/_T_217 ),
        .I4(core_n_0),
        .O(core__161_n_0));
  CARRY4 core__161_i_1
       (.CI(\bypass_mux_1_reg[27]_i_2_n_0 ),
        .CO({core__161_i_1_n_0,core__161_i_1_n_1,core__161_i_1_n_2,core__161_i_1_n_3}),
        .CYINIT(\<const0> ),
        .DI(alu_io_in1[31:28]),
        .O(dcacheArb_io_requestor_1_req_bits_addr[31:28]),
        .S({core__285_n_0,core_rep__12_n_0,core__283_n_0,core__282_n_0}));
  LUT6 #(
    .INIT(64'h0041140014000041)) 
    core__162
       (.I0(core__436_n_0),
        .I1(alu_io_in1[1]),
        .I2(alu_io_in2[1]),
        .I3(ex_ctrl_alu_fn),
        .I4(alu_io_in2[0]),
        .I5(core_n_1782),
        .O(core__162_n_0));
  LUT6 #(
    .INIT(64'h0041140014000041)) 
    core__163
       (.I0(core__439_n_0),
        .I1(alu_io_in1[4]),
        .I2(alu_io_in2[4]),
        .I3(ex_ctrl_alu_fn),
        .I4(alu_io_in2[3]),
        .I5(alu_io_in1[3]),
        .O(core__163_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__164
       (.I0(alu_io_in1[8]),
        .I1(alu_io_in2[8]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[7]),
        .I4(alu_io_in2[7]),
        .I5(core__440_n_0),
        .O(core__164_n_0));
  LUT6 #(
    .INIT(64'h0041140014000041)) 
    core__165
       (.I0(core__441_n_0),
        .I1(alu_io_in1[10]),
        .I2(alu_io_in2[10]),
        .I3(ex_ctrl_alu_fn),
        .I4(alu_io_in2[9]),
        .I5(alu_io_in1[9]),
        .O(core__165_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__166
       (.I0(alu_io_in1[14]),
        .I1(alu_io_in2[14]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[13]),
        .I4(alu_io_in2[13]),
        .I5(core__442_n_0),
        .O(core__166_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__167
       (.I0(alu_io_in1[17]),
        .I1(alu_io_in2[17]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[16]),
        .I4(alu_io_in2[16]),
        .I5(core__443_n_0),
        .O(core__167_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__168
       (.I0(alu_io_in1[20]),
        .I1(alu_io_in2[20]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[19]),
        .I4(alu_io_in2[19]),
        .I5(core__444_n_0),
        .O(core__168_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__169
       (.I0(alu_io_in1[23]),
        .I1(alu_io_in2[23]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[22]),
        .I4(alu_io_in2[22]),
        .I5(core__445_n_0),
        .O(core__169_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__17
       (.I0(_GEN_274[53]),
        .I1(frontend_n_351),
        .I2(_T_1406[53]),
        .I3(frontend_n_352),
        .O(core__17_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__170
       (.I0(alu_io_in1[26]),
        .I1(alu_io_in2[26]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[25]),
        .I4(alu_io_in2[25]),
        .I5(core__446_n_0),
        .O(core__170_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__171
       (.I0(alu_io_in1[29]),
        .I1(alu_io_in2[29]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[28]),
        .I4(alu_io_in2[28]),
        .I5(core__447_n_0),
        .O(core__171_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__172
       (.I0(alu_io_in1[32]),
        .I1(alu_io_in2[32]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[31]),
        .I4(alu_io_in2[31]),
        .I5(core__448_n_0),
        .O(core__172_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__173
       (.I0(alu_io_in1[35]),
        .I1(alu_io_in2[35]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[34]),
        .I4(alu_io_in2[34]),
        .I5(core__449_n_0),
        .O(core__173_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__174
       (.I0(alu_io_in1[38]),
        .I1(alu_io_in2[38]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[37]),
        .I4(alu_io_in2[37]),
        .I5(core__450_n_0),
        .O(core__174_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__175
       (.I0(alu_io_in1[41]),
        .I1(alu_io_in2[41]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[40]),
        .I4(alu_io_in2[40]),
        .I5(core__451_n_0),
        .O(core__175_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__176
       (.I0(alu_io_in1[44]),
        .I1(alu_io_in2[44]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[43]),
        .I4(alu_io_in2[43]),
        .I5(core__452_n_0),
        .O(core__176_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__177
       (.I0(alu_io_in1[47]),
        .I1(alu_io_in2[47]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[46]),
        .I4(alu_io_in2[46]),
        .I5(core__453_n_0),
        .O(core__177_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__178
       (.I0(alu_io_in1[50]),
        .I1(alu_io_in2[50]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[49]),
        .I4(alu_io_in2[49]),
        .I5(core__454_n_0),
        .O(core__178_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__179
       (.I0(alu_io_in1[53]),
        .I1(alu_io_in2[53]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[52]),
        .I4(alu_io_in2[52]),
        .I5(core__455_n_0),
        .O(core__179_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__18
       (.I0(_GEN_274[52]),
        .I1(frontend_n_351),
        .I2(_T_1406[52]),
        .I3(frontend_n_352),
        .O(core__18_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__180
       (.I0(alu_io_in1[56]),
        .I1(alu_io_in2[56]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[55]),
        .I4(alu_io_in2[55]),
        .I5(core__456_n_0),
        .O(core__180_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__181
       (.I0(alu_io_in1[59]),
        .I1(alu_io_in2[59]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[58]),
        .I4(alu_io_in2[58]),
        .I5(core__457_n_0),
        .O(core__181_n_0));
  LUT6 #(
    .INIT(64'h0000000009606009)) 
    core__182
       (.I0(alu_io_in1[62]),
        .I1(alu_io_in2[62]),
        .I2(ex_ctrl_alu_fn),
        .I3(alu_io_in1[61]),
        .I4(alu_io_in2[61]),
        .I5(core__458_n_0),
        .O(core__182_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2478" *) 
  LUT5 #(
    .INIT(32'h00000008)) 
    core__183
       (.I0(ex_ctrl_div),
        .I1(ex_reg_valid),
        .I2(core_n_98),
        .I3(core_n_99),
        .I4(\div/_T_216 ),
        .O(core__183_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2483" *) 
  LUT5 #(
    .INIT(32'hC0FFFFAA)) 
    core__184
       (.I0(\div/_T_216 ),
        .I1(wb_reg_valid),
        .I2(wb_ctrl_wxd),
        .I3(core_n_98),
        .I4(core_n_99),
        .O(core__184_n_0));
  LUT6 #(
    .INIT(64'h0000BA00FFFFFFFF)) 
    core__185
       (.I0(wb_ctrl_div),
        .I1(dcacheArb_io_requestor_1_resp_valid),
        .I2(wb_ctrl_mem),
        .I3(wb_ctrl_wxd),
        .I4(dcache_n_555),
        .I5(core_n_1095),
        .O(core__185_n_0));
  LUT6 #(
    .INIT(64'h01000000FFFFFFFF)) 
    core__186
       (.I0(dcacheArb_io_requestor_1_s2_nack),
        .I1(wb_reg_replay),
        .I2(dcache_io_cpu_invalidate_lr),
        .I3(wb_reg_valid),
        .I4(wb_ctrl_wxd),
        .I5(core_n_1095),
        .O(core__186_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    core__187
       (.I0(core_n_134),
        .I1(\div/_GEN_35 [0]),
        .I2(\div/_GEN_35 [1]),
        .I3(core_n_135),
        .O(core__187_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    core__188
       (.I0(core_n_117),
        .I1(\div/_GEN_35 [0]),
        .I2(core_n_118),
        .I3(\div/_GEN_35 [1]),
        .O(core__188_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    core__189
       (.I0(core_n_168),
        .I1(\div/_GEN_35 [0]),
        .I2(core_n_169),
        .I3(\div/_GEN_35 [1]),
        .O(core__189_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__19
       (.I0(_GEN_274[51]),
        .I1(frontend_n_351),
        .I2(_T_1406[51]),
        .I3(frontend_n_352),
        .O(core__19_n_0));
  LUT4 #(
    .INIT(16'h7888)) 
    core__190
       (.I0(core_n_151),
        .I1(\div/_GEN_35 [0]),
        .I2(core_n_152),
        .I3(\div/_GEN_35 [1]),
        .O(core__190_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2478" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    core__191
       (.I0(core_n_99),
        .I1(core_n_98),
        .I2(\div/_T_216 ),
        .O(core__191_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2483" *) 
  LUT3 #(
    .INIT(8'h04)) 
    core__192
       (.I0(\div/_T_216 ),
        .I1(core_n_99),
        .I2(core_n_98),
        .O(core__192_n_0));
  LUT5 #(
    .INIT(32'h00E2E2E2)) 
    core__193
       (.I0(ex_sfence),
        .I1(core_n_1364),
        .I2(mem_reg_sfence),
        .I3(mem_reg_flush_pipe),
        .I4(mem_reg_valid),
        .O(core__193_n_0));
  LUT5 #(
    .INIT(32'hFCCCAAAA)) 
    core__194
       (.I0(core_n_28),
        .I1(ex_ctrl_fence_i),
        .I2(csr_io_status_debug),
        .I3(ex_ctrl_jalr),
        .I4(mem_ctrl_fp),
        .O(core__194_n_0));
  LUT5 #(
    .INIT(32'hFCCCAAAA)) 
    core__195
       (.I0(mem_reg_flush_pipe),
        .I1(ex_reg_flush_pipe),
        .I2(csr_io_status_debug),
        .I3(ex_ctrl_jalr),
        .I4(mem_ctrl_fp),
        .O(core__195_n_0));
  LUT4 #(
    .INIT(16'hCFAA)) 
    core__196
       (.I0(mem_reg_slow_bypass),
        .I1(core_n_1706),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I3(mem_ctrl_fp),
        .O(core__196_n_0));
  LUT4 #(
    .INIT(16'h4404)) 
    core__197
       (.I0(core_n_1013),
        .I1(core_n_1010),
        .I2(wb_reg_xcpt),
        .I3(wb_reg_cause),
        .O(core__197_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    core__198
       (.I0(wb_reg_xcpt),
        .I1(wb_reg_cause),
        .I2(core_n_1010),
        .I3(core_n_1013),
        .O(core__198_n_0));
  LUT4 #(
    .INIT(16'h0051)) 
    core__199
       (.I0(core_n_1013),
        .I1(wb_reg_xcpt),
        .I2(wb_reg_cause),
        .I3(core_n_1010),
        .O(core__199_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__20
       (.I0(_GEN_274[50]),
        .I1(frontend_n_351),
        .I2(_T_1406[50]),
        .I3(frontend_n_352),
        .O(core__20_n_0));
  LUT4 #(
    .INIT(16'h1FE0)) 
    core__200
       (.I0(mem_ctrl_jal),
        .I1(core_n_1355),
        .I2(_T_20810),
        .I3(mem_reg_pc[32]),
        .O(core__200_n_0));
  LUT6 #(
    .INIT(64'h1110001000000000)) 
    core__201
       (.I0(mem_reg_sfence),
        .I1(csr_io_status_isa[2]),
        .I2(p_0_in[1]),
        .I3(mem_ctrl_jalr),
        .I4(core_n_1331),
        .I5(mem_reg_valid),
        .O(core__201_n_0));
  CARRY4 core__201_i_1
       (.CI(\<const0> ),
        .CO({core__201_i_1_n_0,core__201_i_1_n_1,core__201_i_1_n_2,core__201_i_1_n_3}),
        .CYINIT(\<const0> ),
        .DI({mem_reg_pc[3:1],\<const0> }),
        .O(p_0_in[3:0]),
        .S({core__201_i_2_n_0,core__201_i_3_n_0,core__201_i_4_n_0,\<const0> }));
  LUT5 #(
    .INIT(32'h556AAA6A)) 
    core__201_i_2
       (.I0(mem_reg_pc[3]),
        .I1(core_n_1111),
        .I2(mem_ctrl_jal),
        .I3(core_n_1355),
        .I4(mem_waddr[3]),
        .O(core__201_i_2_n_0));
  LUT6 #(
    .INIT(64'h55556A59AAAA6A59)) 
    core__201_i_3
       (.I0(mem_reg_pc[2]),
        .I1(mem_ctrl_jal),
        .I2(core_n_1112),
        .I3(mem_reg_rvc),
        .I4(core_n_1355),
        .I5(mem_waddr[2]),
        .O(core__201_i_3_n_0));
  LUT6 #(
    .INIT(64'h555556A6AAAA56A6)) 
    core__201_i_4
       (.I0(mem_reg_pc[1]),
        .I1(mem_reg_rvc),
        .I2(mem_ctrl_jal),
        .I3(core_n_1113),
        .I4(core_n_1355),
        .I5(mem_waddr[1]),
        .O(core__201_i_4_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__202
       (.I0(core_n_1557),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__202_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__203
       (.I0(core_n_1556),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__203_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__204
       (.I0(core_n_1555),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__204_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__205
       (.I0(core_n_1554),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__205_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__206
       (.I0(core_n_1553),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__206_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__207
       (.I0(core_n_1552),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__207_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__208
       (.I0(core_n_1551),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__208_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__209
       (.I0(core_n_1550),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__209_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__21
       (.I0(_GEN_274[49]),
        .I1(frontend_n_351),
        .I2(_T_1406[49]),
        .I3(frontend_n_352),
        .O(core__21_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__210
       (.I0(core_n_1549),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__210_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__211
       (.I0(core_n_1548),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__211_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__212
       (.I0(core_n_1547),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__212_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__213
       (.I0(core_n_1546),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__213_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__214
       (.I0(core_n_1545),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__214_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__215
       (.I0(core_n_1544),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__215_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__216
       (.I0(core_n_1543),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__216_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__217
       (.I0(core_n_1542),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__217_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__218
       (.I0(core_n_1541),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__218_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__219
       (.I0(core_n_1540),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__219_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__22
       (.I0(_GEN_274[48]),
        .I1(frontend_n_351),
        .I2(_T_1406[48]),
        .I3(frontend_n_352),
        .O(core__22_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__220
       (.I0(core_n_1539),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__220_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__221
       (.I0(core_n_1538),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__221_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__222
       (.I0(core_n_1537),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__222_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__223
       (.I0(core_n_1536),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__223_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__224
       (.I0(core_n_1535),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__224_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__225
       (.I0(core_n_1534),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__225_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__226
       (.I0(core_n_1533),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__226_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__227
       (.I0(core_n_1532),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__227_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__228
       (.I0(core_n_1531),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__228_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__229
       (.I0(core_n_1530),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__229_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__23
       (.I0(_GEN_274[47]),
        .I1(frontend_n_351),
        .I2(_T_1406[47]),
        .I3(frontend_n_352),
        .O(core__23_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__230
       (.I0(core_n_1529),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__230_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__231
       (.I0(core_n_1528),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__231_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__232
       (.I0(core_n_1527),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__232_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__233
       (.I0(core_n_1526),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__233_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__234
       (.I0(core_n_1525),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__234_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__235
       (.I0(core_n_1524),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__235_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__236
       (.I0(core_n_1523),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__236_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__237
       (.I0(core_n_1522),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__237_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__238
       (.I0(core_n_1521),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__238_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__239
       (.I0(core_n_1520),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__239_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__24
       (.I0(_GEN_274[46]),
        .I1(frontend_n_351),
        .I2(_T_1406[46]),
        .I3(frontend_n_352),
        .O(core__24_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__240
       (.I0(core_n_1519),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__240_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__241
       (.I0(core_n_1518),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__241_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__242
       (.I0(core_n_1517),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__242_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__243
       (.I0(core_n_1516),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__243_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__244
       (.I0(core_n_1515),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__244_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__245
       (.I0(core_n_1514),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__245_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__246
       (.I0(core_n_1513),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__246_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__247
       (.I0(core_n_1512),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__247_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__248
       (.I0(core_n_1511),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__248_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__249
       (.I0(core_n_1510),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__249_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__25
       (.I0(_GEN_274[45]),
        .I1(frontend_n_351),
        .I2(_T_1406[45]),
        .I3(frontend_n_352),
        .O(core__25_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__250
       (.I0(core_n_1509),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__250_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__251
       (.I0(core_n_1508),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__251_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__252
       (.I0(core_n_1507),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__252_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__253
       (.I0(core_n_1506),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__253_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__254
       (.I0(core_n_1505),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__254_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__255
       (.I0(core_n_1504),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__255_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__256
       (.I0(core_n_1503),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__256_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__257
       (.I0(core_n_1502),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__257_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__258
       (.I0(core_n_1501),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__258_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__259
       (.I0(core_n_1500),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__259_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__26
       (.I0(_GEN_274[44]),
        .I1(frontend_n_351),
        .I2(_T_1406[44]),
        .I3(frontend_n_352),
        .O(core__26_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__260
       (.I0(core_n_1499),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__260_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__261
       (.I0(core_n_1498),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__261_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__262
       (.I0(core_n_1497),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__262_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__263
       (.I0(core_n_1496),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__263_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core__264
       (.I0(core_n_1495),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core__264_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2484" *) 
  LUT3 #(
    .INIT(8'h04)) 
    core__265
       (.I0(core_n_1346),
        .I1(core_n_1345),
        .I2(core_n_1347),
        .O(core__265_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8FFFFFF)) 
    core__266
       (.I0(_T_1944),
        .I1(core_n_30),
        .I2(core_n_1349),
        .I3(core_n_1346),
        .I4(core_n_1345),
        .I5(core_n_1347),
        .O(core__266_n_0));
  CARRY4 core__266_i_1
       (.CI(core__266_i_3_n_0),
        .CO({_T_1944,core__266_i_1_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,core__266_i_4_n_0,core_n_1607}));
  CARRY4 core__266_i_11
       (.CI(core__266_i_16_n_0),
        .CO({core__266_i_11_n_0,core__266_i_11_n_1,core__266_i_11_n_2,core__266_i_11_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1595,core_n_1596,core_n_1597,core_n_1598}));
  CARRY4 core__266_i_16
       (.CI(core__266_i_21_n_0),
        .CO({core__266_i_16_n_0,core__266_i_16_n_1,core__266_i_16_n_2,core__266_i_16_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1591,core_n_1592,core_n_1593,core_n_1594}));
  CARRY4 core__266_i_21
       (.CI(\<const0> ),
        .CO({core__266_i_21_n_0,core__266_i_21_n_1,core__266_i_21_n_2,core__266_i_21_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1490,core_n_1491,core_n_1492,core_n_1493}));
  CARRY4 core__266_i_3
       (.CI(core__266_i_6_n_0),
        .CO({core__266_i_3_n_0,core__266_i_3_n_1,core__266_i_3_n_2,core__266_i_3_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1603,core_n_1604,core_n_1605,core_n_1606}));
  LUT1 #(
    .INIT(2'h1)) 
    core__266_i_4
       (.I0(core_n_1494),
        .O(core__266_i_4_n_0));
  CARRY4 core__266_i_6
       (.CI(core__266_i_11_n_0),
        .CO({core__266_i_6_n_0,core__266_i_6_n_1,core__266_i_6_n_2,core__266_i_6_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1599,core_n_1600,core_n_1601,core_n_1602}));
  LUT3 #(
    .INIT(8'h96)) 
    core__267
       (.I0(alu_io_in1[41]),
        .I1(alu_io_in2[41]),
        .I2(ex_ctrl_alu_fn),
        .O(core__267_n_0));
  LUT6 #(
    .INIT(64'h65AA65659A559A9A)) 
    core__268
       (.I0(alu_io_in1[7]),
        .I1(core_n_1777),
        .I2(mem_reg_rs2[7]),
        .I3(core_n_1776),
        .I4(core_n_1242),
        .I5(ex_ctrl_alu_fn),
        .O(core__268_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__269
       (.I0(alu_io_in1[8]),
        .I1(alu_io_in2[8]),
        .I2(ex_ctrl_alu_fn),
        .O(core__269_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__27
       (.I0(_GEN_274[43]),
        .I1(frontend_n_351),
        .I2(_T_1406[43]),
        .I3(frontend_n_352),
        .O(core__27_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__270
       (.I0(alu_io_in1[9]),
        .I1(alu_io_in2[9]),
        .I2(ex_ctrl_alu_fn),
        .O(core__270_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__271
       (.I0(alu_io_in1[10]),
        .I1(alu_io_in2[10]),
        .I2(ex_ctrl_alu_fn),
        .O(core__271_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__272
       (.I0(alu_io_in1[13]),
        .I1(alu_io_in2[13]),
        .I2(ex_ctrl_alu_fn),
        .O(core__272_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__273
       (.I0(alu_io_in1[14]),
        .I1(alu_io_in2[14]),
        .I2(ex_ctrl_alu_fn),
        .O(core__273_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__274
       (.I0(alu_io_in1[16]),
        .I1(alu_io_in2[16]),
        .I2(ex_ctrl_alu_fn),
        .O(core__274_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__275
       (.I0(alu_io_in1[17]),
        .I1(alu_io_in2[17]),
        .I2(ex_ctrl_alu_fn),
        .O(core__275_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__276
       (.I0(alu_io_in1[19]),
        .I1(alu_io_in2[19]),
        .I2(ex_ctrl_alu_fn),
        .O(core__276_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__277
       (.I0(alu_io_in1[20]),
        .I1(alu_io_in2[20]),
        .I2(ex_ctrl_alu_fn),
        .O(core__277_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__278
       (.I0(alu_io_in1[22]),
        .I1(alu_io_in2[22]),
        .I2(ex_ctrl_alu_fn),
        .O(core__278_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__279
       (.I0(alu_io_in1[23]),
        .I1(alu_io_in2[23]),
        .I2(ex_ctrl_alu_fn),
        .O(core__279_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__28
       (.I0(_GEN_274[42]),
        .I1(frontend_n_351),
        .I2(_T_1406[42]),
        .I3(frontend_n_352),
        .O(core__28_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__280
       (.I0(alu_io_in1[25]),
        .I1(alu_io_in2[25]),
        .I2(ex_ctrl_alu_fn),
        .O(core__280_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__281
       (.I0(alu_io_in1[26]),
        .I1(alu_io_in2[26]),
        .I2(ex_ctrl_alu_fn),
        .O(core__281_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__282
       (.I0(alu_io_in1[28]),
        .I1(alu_io_in2[28]),
        .I2(ex_ctrl_alu_fn),
        .O(core__282_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__283
       (.I0(alu_io_in1[29]),
        .I1(alu_io_in2[29]),
        .I2(ex_ctrl_alu_fn),
        .O(core__283_n_0));
  LUT5 #(
    .INIT(32'h0A800080)) 
    core__284
       (.I0(ex_ctrl_alu_fn),
        .I1(ex_reg_pc),
        .I2(core_n_1680),
        .I3(core_n_1681),
        .I4(core_n_237),
        .O(core__284_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__285
       (.I0(alu_io_in1[31]),
        .I1(alu_io_in2[31]),
        .I2(ex_ctrl_alu_fn),
        .O(core__285_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__286
       (.I0(alu_io_in1[32]),
        .I1(alu_io_in2[32]),
        .I2(ex_ctrl_alu_fn),
        .O(core__286_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__287
       (.I0(alu_io_in1[34]),
        .I1(alu_io_in2[34]),
        .I2(ex_ctrl_alu_fn),
        .O(core__287_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__288
       (.I0(alu_io_in1[35]),
        .I1(alu_io_in2[35]),
        .I2(ex_ctrl_alu_fn),
        .O(core__288_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__289
       (.I0(alu_io_in1[37]),
        .I1(alu_io_in2[37]),
        .I2(ex_ctrl_alu_fn),
        .O(core__289_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__29
       (.I0(_GEN_274[41]),
        .I1(frontend_n_351),
        .I2(_T_1406[41]),
        .I3(frontend_n_352),
        .O(core__29_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__290
       (.I0(alu_io_in1[38]),
        .I1(alu_io_in2[38]),
        .I2(ex_ctrl_alu_fn),
        .O(core__290_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2496" *) 
  LUT2 #(
    .INIT(4'h2)) 
    core__291
       (.I0(core_n_0),
        .I1(core_n_289),
        .O(core__291_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__292
       (.I0(alu_io_in1[63]),
        .I1(alu_io_in2[63]),
        .I2(ex_ctrl_alu_fn),
        .O(core__292_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__293
       (.I0(alu_io_in1[61]),
        .I1(alu_io_in2[61]),
        .I2(ex_ctrl_alu_fn),
        .O(core__293_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__294
       (.I0(alu_io_in1[62]),
        .I1(alu_io_in2[62]),
        .I2(ex_ctrl_alu_fn),
        .O(core__294_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__295
       (.I0(alu_io_in1[58]),
        .I1(alu_io_in2[58]),
        .I2(ex_ctrl_alu_fn),
        .O(core__295_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__296
       (.I0(alu_io_in1[59]),
        .I1(alu_io_in2[59]),
        .I2(ex_ctrl_alu_fn),
        .O(core__296_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__297
       (.I0(alu_io_in1[55]),
        .I1(alu_io_in2[55]),
        .I2(ex_ctrl_alu_fn),
        .O(core__297_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__298
       (.I0(alu_io_in1[56]),
        .I1(alu_io_in2[56]),
        .I2(ex_ctrl_alu_fn),
        .O(core__298_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__299
       (.I0(alu_io_in1[52]),
        .I1(alu_io_in2[52]),
        .I2(ex_ctrl_alu_fn),
        .O(core__299_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__30
       (.I0(_GEN_274[40]),
        .I1(frontend_n_351),
        .I2(_T_1406[40]),
        .I3(frontend_n_352),
        .O(core__30_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__300
       (.I0(alu_io_in1[53]),
        .I1(alu_io_in2[53]),
        .I2(ex_ctrl_alu_fn),
        .O(core__300_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__301
       (.I0(alu_io_in1[49]),
        .I1(alu_io_in2[49]),
        .I2(ex_ctrl_alu_fn),
        .O(core__301_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__302
       (.I0(alu_io_in1[50]),
        .I1(alu_io_in2[50]),
        .I2(ex_ctrl_alu_fn),
        .O(core__302_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__303
       (.I0(alu_io_in1[46]),
        .I1(alu_io_in2[46]),
        .I2(ex_ctrl_alu_fn),
        .O(core__303_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__304
       (.I0(alu_io_in1[47]),
        .I1(alu_io_in2[47]),
        .I2(ex_ctrl_alu_fn),
        .O(core__304_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__305
       (.I0(alu_io_in1[43]),
        .I1(alu_io_in2[43]),
        .I2(ex_ctrl_alu_fn),
        .O(core__305_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__306
       (.I0(alu_io_in1[44]),
        .I1(alu_io_in2[44]),
        .I2(ex_ctrl_alu_fn),
        .O(core__306_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__307
       (.I0(alu_io_in1[40]),
        .I1(alu_io_in2[40]),
        .I2(ex_ctrl_alu_fn),
        .O(core__307_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    core__308
       (.I0(_T_2518[0]),
        .I1(_T_2518[1]),
        .I2(_T_2518[2]),
        .O(core__308_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    core__309
       (.I0(_T_2518[3]),
        .I1(_T_2518[4]),
        .I2(_T_2518[5]),
        .O(core__309_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__31
       (.I0(_GEN_274[39]),
        .I1(frontend_n_351),
        .I2(_T_1406[39]),
        .I3(frontend_n_352),
        .O(core__31_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    core__310
       (.I0(_T_2518[6]),
        .I1(_T_2518[7]),
        .I2(_T_2518[8]),
        .O(core__310_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    core__311
       (.I0(_T_2518[9]),
        .I1(_T_2518[10]),
        .I2(_T_2518[11]),
        .O(core__311_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    core__312
       (.I0(_T_2518[12]),
        .I1(_T_2518[13]),
        .I2(_T_2518[14]),
        .O(core__312_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    core__313
       (.I0(_T_2518[15]),
        .I1(_T_2518[16]),
        .I2(_T_2518[17]),
        .O(core__313_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    core__314
       (.I0(_T_2518[18]),
        .I1(_T_2518[19]),
        .I2(_T_2518[20]),
        .O(core__314_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    core__315
       (.I0(_T_2518[21]),
        .I1(_T_2518[22]),
        .I2(_T_2518[23]),
        .O(core__315_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2559" *) 
  LUT3 #(
    .INIT(8'h40)) 
    core__316
       (.I0(wb_waddr[2]),
        .I1(wb_waddr[1]),
        .I2(wb_waddr[0]),
        .O(core__316_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2560" *) 
  LUT3 #(
    .INIT(8'h04)) 
    core__317
       (.I0(wb_waddr[2]),
        .I1(wb_waddr[1]),
        .I2(wb_waddr[0]),
        .O(core__317_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2559" *) 
  LUT3 #(
    .INIT(8'h04)) 
    core__318
       (.I0(wb_waddr[2]),
        .I1(wb_waddr[0]),
        .I2(wb_waddr[1]),
        .O(core__318_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2560" *) 
  LUT3 #(
    .INIT(8'h01)) 
    core__319
       (.I0(wb_waddr[2]),
        .I1(wb_waddr[1]),
        .I2(wb_waddr[0]),
        .O(core__319_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__32
       (.I0(_GEN_274[38]),
        .I1(frontend_n_351),
        .I2(_T_1406[38]),
        .I3(frontend_n_352),
        .O(core__32_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__320
       (.I0(ex_ctrl_alu_fn),
        .I1(alu_io_in2[0]),
        .O(core__320_n_0));
  LUT6 #(
    .INIT(64'hBF00000000000000)) 
    core__321
       (.I0(ex_ctrl_sel_imm[1]),
        .I1(ex_ctrl_sel_imm[2]),
        .I2(ex_ctrl_sel_imm[0]),
        .I3(_T_1686),
        .I4(ex_ctrl_sel_alu2[0]),
        .I5(ex_ctrl_sel_alu2[1]),
        .O(core__321_n_0));
  LUT3 #(
    .INIT(8'h40)) 
    core__322
       (.I0(ex_ctrl_sel_imm[1]),
        .I1(ex_ctrl_sel_imm[2]),
        .I2(ex_ctrl_sel_imm[0]),
        .O(core__322_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    core__323
       (.I0(core_n_1329),
        .I1(csr_io_bp_0_address[38]),
        .O(core__323_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__324
       (.I0(\div/_GEN_36 [63]),
        .I1(core_n_105),
        .O(core__324_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__325
       (.I0(core_n_357),
        .I1(core_n_371),
        .O(core__325_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__326
       (.I0(core_n_357),
        .I1(core_n_372),
        .O(core__326_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__327
       (.I0(core_n_357),
        .I1(core_n_373),
        .O(core__327_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__328
       (.I0(core_n_357),
        .I1(core_n_366),
        .O(core__328_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__329
       (.I0(core_n_357),
        .I1(core_n_367),
        .O(core__329_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__33
       (.I0(_GEN_274[37]),
        .I1(frontend_n_351),
        .I2(_T_1406[37]),
        .I3(frontend_n_352),
        .O(core__33_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__330
       (.I0(core_n_357),
        .I1(core_n_368),
        .O(core__330_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__331
       (.I0(core_n_357),
        .I1(core_n_369),
        .O(core__331_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__332
       (.I0(core_n_357),
        .I1(core_n_362),
        .O(core__332_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__333
       (.I0(core_n_357),
        .I1(core_n_363),
        .O(core__333_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__334
       (.I0(core_n_357),
        .I1(core_n_364),
        .O(core__334_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__335
       (.I0(core_n_357),
        .I1(core_n_365),
        .O(core__335_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__336
       (.I0(core_n_357),
        .I1(core_n_358),
        .O(core__336_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__337
       (.I0(core_n_357),
        .I1(core_n_359),
        .O(core__337_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__338
       (.I0(core_n_357),
        .I1(core_n_360),
        .O(core__338_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__339
       (.I0(core_n_357),
        .I1(core_n_361),
        .O(core__339_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__34
       (.I0(_GEN_274[36]),
        .I1(frontend_n_351),
        .I2(_T_1406[36]),
        .I3(frontend_n_352),
        .O(core__34_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__340
       (.I0(core_n_357),
        .I1(core_n_375),
        .O(core__340_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__341
       (.I0(core_n_357),
        .I1(core_n_370),
        .O(core__341_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__342
       (.I0(core_n_387),
        .I1(core_n_356),
        .O(core__342_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__342_i_10
       (.I0(core_n_327),
        .I1(core_n_336),
        .O(core__342_i_10_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    core__342_i_12
       (.I0(core_n_357),
        .O(core__342_i_12_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    core__342_i_13
       (.I0(core_n_357),
        .O(core__342_i_13_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    core__342_i_14
       (.I0(core_n_357),
        .O(core__342_i_14_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    core__342_i_15
       (.I0(core_n_357),
        .O(core__342_i_15_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    core__342_i_20
       (.I0(core_n_357),
        .O(core__342_i_20_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    core__342_i_21
       (.I0(core_n_357),
        .O(core__342_i_21_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    core__342_i_22
       (.I0(core_n_357),
        .O(core__342_i_22_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    core__342_i_23
       (.I0(core_n_357),
        .O(core__342_i_23_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    core__342_i_4
       (.I0(core_n_357),
        .O(core__342_i_4_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    core__342_i_5
       (.I0(core_n_357),
        .O(core__342_i_5_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__342_i_6
       (.I0(core_n_374),
        .I1(core_n_357),
        .O(core__342_i_6_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__342_i_8
       (.I0(core_n_327),
        .I1(core_n_340),
        .O(core__342_i_8_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__342_i_9
       (.I0(core_n_327),
        .I1(core_n_341),
        .O(core__342_i_9_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__343
       (.I0(core_n_387),
        .I1(core_n_350),
        .O(core__343_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__343_i_2
       (.I0(core_n_327),
        .I1(core_n_337),
        .O(core__343_i_2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__343_i_3
       (.I0(core_n_327),
        .I1(core_n_338),
        .O(core__343_i_3_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__343_i_4
       (.I0(core_n_327),
        .I1(core_n_339),
        .O(core__343_i_4_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__343_i_5
       (.I0(core_n_327),
        .I1(core_n_332),
        .O(core__343_i_5_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__344
       (.I0(core_n_387),
        .I1(core_n_351),
        .O(core__344_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__345
       (.I0(core_n_387),
        .I1(core_n_352),
        .O(core__345_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__346
       (.I0(core_n_387),
        .I1(core_n_353),
        .O(core__346_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__347
       (.I0(core_n_387),
        .I1(core_n_346),
        .O(core__347_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__347_i_2
       (.I0(core_n_327),
        .I1(core_n_333),
        .O(core__347_i_2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__347_i_3
       (.I0(core_n_327),
        .I1(core_n_334),
        .O(core__347_i_3_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__347_i_4
       (.I0(core_n_327),
        .I1(core_n_335),
        .O(core__347_i_4_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__347_i_5
       (.I0(core_n_327),
        .I1(core_n_328),
        .O(core__347_i_5_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__348
       (.I0(core_n_387),
        .I1(core_n_347),
        .O(core__348_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__349
       (.I0(core_n_387),
        .I1(core_n_348),
        .O(core__349_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__35
       (.I0(_GEN_274[35]),
        .I1(frontend_n_351),
        .I2(_T_1406[35]),
        .I3(frontend_n_352),
        .O(core__35_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__350
       (.I0(core_n_387),
        .I1(core_n_349),
        .O(core__350_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__351
       (.I0(core_n_387),
        .I1(core_n_342),
        .O(core__351_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__351_i_2
       (.I0(core_n_327),
        .I1(core_n_329),
        .O(core__351_i_2_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__351_i_3
       (.I0(core_n_327),
        .I1(core_n_330),
        .O(core__351_i_3_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__351_i_4
       (.I0(core_n_327),
        .I1(core_n_331),
        .O(core__351_i_4_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__352
       (.I0(core_n_387),
        .I1(core_n_343),
        .O(core__352_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__353
       (.I0(core_n_387),
        .I1(core_n_344),
        .O(core__353_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__354
       (.I0(core_n_387),
        .I1(core_n_345),
        .O(core__354_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__355
       (.I0(core_n_387),
        .I1(core_n_323),
        .O(core__355_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__356
       (.I0(core_n_387),
        .I1(core_n_324),
        .O(core__356_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__357
       (.I0(core_n_387),
        .I1(core_n_325),
        .O(core__357_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__358
       (.I0(O),
        .I1(core_n_354),
        .O(core__358_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__359
       (.I0(O),
        .I1(core_n_387),
        .O(core__359_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__36
       (.I0(_GEN_274[34]),
        .I1(frontend_n_351),
        .I2(_T_1406[34]),
        .I3(frontend_n_352),
        .O(core__36_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__360
       (.I0(\div/_GEN_36 [62]),
        .I1(\div/_T_103 ),
        .O(core__360_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__361
       (.I0(\div/_GEN_36 [61]),
        .I1(core_n_107),
        .O(core__361_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__362
       (.I0(\div/_GEN_36 [60]),
        .I1(core_n_108),
        .O(core__362_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__363
       (.I0(\div/_GEN_36 [59]),
        .I1(core_n_109),
        .O(core__363_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__364
       (.I0(\div/_GEN_36 [58]),
        .I1(core_n_110),
        .O(core__364_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__365
       (.I0(\div/_GEN_36 [57]),
        .I1(core_n_111),
        .O(core__365_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__366
       (.I0(\div/_GEN_36 [56]),
        .I1(core_n_112),
        .O(core__366_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__367
       (.I0(\div/_GEN_36 [55]),
        .I1(core_n_113),
        .O(core__367_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__368
       (.I0(\div/_GEN_36 [54]),
        .I1(core_n_114),
        .O(core__368_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__369
       (.I0(\div/_GEN_36 [53]),
        .I1(core_n_115),
        .O(core__369_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__37
       (.I0(_GEN_274[33]),
        .I1(frontend_n_351),
        .I2(_T_1406[33]),
        .I3(frontend_n_352),
        .O(core__37_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__370
       (.I0(\div/_GEN_36 [52]),
        .I1(core_n_116),
        .O(core__370_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__371
       (.I0(\div/_GEN_36 [51]),
        .I1(core_n_117),
        .O(core__371_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__372
       (.I0(\div/_GEN_36 [50]),
        .I1(core_n_118),
        .O(core__372_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__373
       (.I0(\div/_GEN_36 [49]),
        .I1(core_n_119),
        .O(core__373_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__374
       (.I0(\div/_GEN_36 [48]),
        .I1(core_n_120),
        .O(core__374_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__375
       (.I0(\div/_GEN_36 [47]),
        .I1(core_n_121),
        .O(core__375_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__376
       (.I0(\div/_GEN_36 [46]),
        .I1(core_n_122),
        .O(core__376_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__377
       (.I0(\div/_GEN_36 [45]),
        .I1(core_n_123),
        .O(core__377_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__378
       (.I0(\div/_GEN_36 [44]),
        .I1(core_n_124),
        .O(core__378_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__379
       (.I0(\div/_GEN_36 [43]),
        .I1(core_n_125),
        .O(core__379_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__38
       (.I0(_GEN_274[32]),
        .I1(frontend_n_351),
        .I2(_T_1406[32]),
        .I3(frontend_n_352),
        .O(core__38_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__380
       (.I0(\div/_GEN_36 [42]),
        .I1(core_n_126),
        .O(core__380_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__381
       (.I0(\div/_GEN_36 [41]),
        .I1(core_n_127),
        .O(core__381_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__382
       (.I0(\div/_GEN_36 [40]),
        .I1(core_n_128),
        .O(core__382_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__383
       (.I0(\div/_GEN_36 [39]),
        .I1(core_n_129),
        .O(core__383_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__384
       (.I0(\div/_GEN_36 [38]),
        .I1(core_n_130),
        .O(core__384_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__385
       (.I0(\div/_GEN_36 [37]),
        .I1(core_n_131),
        .O(core__385_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__386
       (.I0(\div/_GEN_36 [36]),
        .I1(core_n_132),
        .O(core__386_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__387
       (.I0(\div/_GEN_36 [35]),
        .I1(core_n_133),
        .O(core__387_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__388
       (.I0(\div/_GEN_36 [34]),
        .I1(core_n_134),
        .O(core__388_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__389
       (.I0(\div/_GEN_36 [33]),
        .I1(core_n_135),
        .O(core__389_n_0));
  LUT5 #(
    .INIT(32'h55545555)) 
    core__39
       (.I0(_T_1142[13]),
        .I1(frontend_n_370),
        .I2(frontend_n_369),
        .I3(frontend_n_368),
        .I4(frontend_n_371),
        .O(core__39_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__390
       (.I0(\div/_GEN_36 [32]),
        .I1(core_n_136),
        .O(core__390_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__391
       (.I0(\div/_GEN_36 [31]),
        .I1(core_n_137),
        .O(core__391_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__392
       (.I0(\div/_GEN_36 [30]),
        .I1(core_n_138),
        .O(core__392_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__393
       (.I0(\div/_GEN_36 [29]),
        .I1(core_n_139),
        .O(core__393_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__394
       (.I0(\div/_GEN_36 [28]),
        .I1(core_n_140),
        .O(core__394_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__395
       (.I0(\div/_GEN_36 [27]),
        .I1(core_n_141),
        .O(core__395_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__396
       (.I0(\div/_GEN_36 [26]),
        .I1(core_n_142),
        .O(core__396_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__397
       (.I0(\div/_GEN_36 [25]),
        .I1(core_n_143),
        .O(core__397_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__398
       (.I0(\div/_GEN_36 [24]),
        .I1(core_n_144),
        .O(core__398_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__399
       (.I0(\div/_GEN_36 [23]),
        .I1(core_n_145),
        .O(core__399_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2499" *) 
  LUT4 #(
    .INIT(16'hC0AA)) 
    core__4
       (.I0(core_n_32),
        .I1(_T_1829),
        .I2(frontend_n_352),
        .I3(_T_1790),
        .O(core__4_n_0));
  LUT6 #(
    .INIT(64'h0000000001010001)) 
    core__40
       (.I0(frontend_n_396),
        .I1(_T_1005[6]),
        .I2(_T_1050[2]),
        .I3(_T_1142[30]),
        .I4(_T_1031[14]),
        .I5(id_ctrl_alu_dw),
        .O(core__40_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__400
       (.I0(\div/_GEN_36 [22]),
        .I1(core_n_146),
        .O(core__400_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__401
       (.I0(\div/_GEN_36 [21]),
        .I1(core_n_147),
        .O(core__401_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__402
       (.I0(\div/_GEN_36 [20]),
        .I1(core_n_148),
        .O(core__402_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__403
       (.I0(\div/_GEN_36 [19]),
        .I1(core_n_149),
        .O(core__403_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__404
       (.I0(\div/_GEN_36 [18]),
        .I1(core_n_150),
        .O(core__404_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__405
       (.I0(\div/_GEN_36 [17]),
        .I1(core_n_151),
        .O(core__405_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__406
       (.I0(\div/_GEN_36 [16]),
        .I1(core_n_152),
        .O(core__406_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__407
       (.I0(\div/_GEN_36 [15]),
        .I1(core_n_153),
        .O(core__407_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__408
       (.I0(\div/_GEN_36 [14]),
        .I1(core_n_154),
        .O(core__408_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__409
       (.I0(\div/_GEN_36 [13]),
        .I1(core_n_155),
        .O(core__409_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2544" *) 
  LUT3 #(
    .INIT(8'h15)) 
    core__41
       (.I0(_T_1142[13]),
        .I1(_T_1142[30]),
        .I2(_T_1142[12]),
        .O(core__41_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__410
       (.I0(\div/_GEN_36 [12]),
        .I1(core_n_156),
        .O(core__410_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__411
       (.I0(\div/_GEN_36 [11]),
        .I1(core_n_157),
        .O(core__411_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__412
       (.I0(\div/_GEN_36 [10]),
        .I1(core_n_158),
        .O(core__412_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__413
       (.I0(\div/_GEN_36 [9]),
        .I1(core_n_159),
        .O(core__413_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__414
       (.I0(\div/_GEN_36 [8]),
        .I1(core_n_160),
        .O(core__414_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__415
       (.I0(\div/_GEN_36 [7]),
        .I1(core_n_161),
        .O(core__415_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__416
       (.I0(\div/_GEN_36 [6]),
        .I1(core_n_162),
        .O(core__416_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__417
       (.I0(\div/_GEN_36 [5]),
        .I1(core_n_163),
        .O(core__417_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__418
       (.I0(\div/_GEN_36 [4]),
        .I1(core_n_164),
        .O(core__418_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__419
       (.I0(\div/_GEN_36 [3]),
        .I1(core_n_165),
        .O(core__419_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    core__42
       (.I0(frontend_n_378),
        .I1(frontend_n_396),
        .O(core__42_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__420
       (.I0(\div/_GEN_36 [2]),
        .I1(core_n_166),
        .O(core__420_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__421
       (.I0(\div/_GEN_36 [1]),
        .I1(core_n_167),
        .O(core__421_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__422
       (.I0(\div/_GEN_36 [0]),
        .I1(core_n_168),
        .O(core__422_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__423
       (.I0(\div/_GEN_35 [1]),
        .I1(core_n_169),
        .O(core__423_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__424
       (.I0(mem_reg_pc[32]),
        .I1(mem_reg_pc[33]),
        .O(core__424_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__425
       (.I0(mem_reg_pc[33]),
        .I1(mem_reg_pc[34]),
        .O(core__425_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__426
       (.I0(mem_reg_pc[34]),
        .I1(mem_reg_pc[35]),
        .O(core__426_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__427
       (.I0(mem_reg_pc[35]),
        .I1(mem_reg_pc[36]),
        .O(core__427_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__428
       (.I0(mem_reg_pc[36]),
        .I1(mem_reg_pc[37]),
        .O(core__428_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__429
       (.I0(mem_reg_pc[38]),
        .I1(mem_reg_pc[39]),
        .O(core__429_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    core__43
       (.I0(_T_1031[14]),
        .I1(_T_1050[5]),
        .O(core__43_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__430
       (.I0(mem_reg_pc[37]),
        .I1(mem_reg_pc[38]),
        .O(core__430_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__431
       (.I0(_GEN_277[62]),
        .I1(dcacheArb_io_requestor_1_s1_data_data[63]),
        .O(core__431_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__432
       (.I0(_GEN_277[126]),
        .I1(dcacheArb_io_requestor_1_s1_data_data[63]),
        .O(core__432_n_0));
  LUT5 #(
    .INIT(32'hBBBBBBB0)) 
    core__433
       (.I0(wb_reg_cause),
        .I1(wb_reg_xcpt),
        .I2(core__121_n_0),
        .I3(csr_io_rw_addr[1]),
        .I4(csr_io_rw_addr[2]),
        .O(core__433_n_0));
  LUT4 #(
    .INIT(16'hF444)) 
    core__434
       (.I0(core_n_1350),
        .I1(core_n_30),
        .I2(core_n_1365),
        .I3(core_n_1349),
        .O(core__434_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core__435
       (.I0(alu_io_in1[1]),
        .I1(alu_io_in2[1]),
        .I2(ex_ctrl_alu_fn),
        .O(core__435_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2543" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__436
       (.I0(alu_io_in1[2]),
        .I1(alu_io_in2[2]),
        .I2(ex_ctrl_alu_fn),
        .O(core__436_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2558" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__437
       (.I0(alu_io_in1[3]),
        .I1(alu_io_in2[3]),
        .I2(ex_ctrl_alu_fn),
        .O(core__437_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2558" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__438
       (.I0(alu_io_in1[4]),
        .I1(alu_io_in2[4]),
        .I2(ex_ctrl_alu_fn),
        .O(core__438_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2550" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__439
       (.I0(alu_io_in1[5]),
        .I1(alu_io_in2[5]),
        .I2(ex_ctrl_alu_fn),
        .O(core__439_n_0));
  LUT6 #(
    .INIT(64'h5555555545405555)) 
    core__44
       (.I0(frontend_n_232),
        .I1(_T_1406[0]),
        .I2(frontend_n_351),
        .I3(_GEN_274[0]),
        .I4(frontend_n_388),
        .I5(_T_1829),
        .O(core__44_n_0));
  LUT6 #(
    .INIT(64'h65AA65659A559A9A)) 
    core__440
       (.I0(alu_io_in1[6]),
        .I1(core_n_1777),
        .I2(mem_reg_rs2[6]),
        .I3(core_n_1776),
        .I4(core_n_1243),
        .I5(ex_ctrl_alu_fn),
        .O(core__440_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2555" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__441
       (.I0(alu_io_in1[11]),
        .I1(alu_io_in2[11]),
        .I2(ex_ctrl_alu_fn),
        .O(core__441_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2554" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__442
       (.I0(alu_io_in1[12]),
        .I1(alu_io_in2[12]),
        .I2(ex_ctrl_alu_fn),
        .O(core__442_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2552" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__443
       (.I0(alu_io_in1[15]),
        .I1(alu_io_in2[15]),
        .I2(ex_ctrl_alu_fn),
        .O(core__443_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2557" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__444
       (.I0(alu_io_in1[18]),
        .I1(alu_io_in2[18]),
        .I2(ex_ctrl_alu_fn),
        .O(core__444_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2557" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__445
       (.I0(alu_io_in1[21]),
        .I1(alu_io_in2[21]),
        .I2(ex_ctrl_alu_fn),
        .O(core__445_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2555" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__446
       (.I0(alu_io_in1[24]),
        .I1(alu_io_in2[24]),
        .I2(ex_ctrl_alu_fn),
        .O(core__446_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2554" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__447
       (.I0(alu_io_in1[27]),
        .I1(alu_io_in2[27]),
        .I2(ex_ctrl_alu_fn),
        .O(core__447_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2550" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__448
       (.I0(alu_io_in1[30]),
        .I1(alu_io_in2[30]),
        .I2(ex_ctrl_alu_fn),
        .O(core__448_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2546" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__449
       (.I0(alu_io_in1[33]),
        .I1(alu_io_in2[33]),
        .I2(ex_ctrl_alu_fn),
        .O(core__449_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2495" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    core__45
       (.I0(_T_1142[12]),
        .I1(_T_1142[13]),
        .I2(_T_1031[14]),
        .I3(_T_1005[6]),
        .O(core__45_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2547" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__450
       (.I0(alu_io_in1[36]),
        .I1(alu_io_in2[36]),
        .I2(ex_ctrl_alu_fn),
        .O(core__450_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2546" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__451
       (.I0(alu_io_in1[39]),
        .I1(alu_io_in2[39]),
        .I2(ex_ctrl_alu_fn),
        .O(core__451_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2549" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__452
       (.I0(alu_io_in1[42]),
        .I1(alu_io_in2[42]),
        .I2(ex_ctrl_alu_fn),
        .O(core__452_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2549" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__453
       (.I0(alu_io_in1[45]),
        .I1(alu_io_in2[45]),
        .I2(ex_ctrl_alu_fn),
        .O(core__453_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2548" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__454
       (.I0(alu_io_in1[48]),
        .I1(alu_io_in2[48]),
        .I2(ex_ctrl_alu_fn),
        .O(core__454_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2548" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__455
       (.I0(alu_io_in1[51]),
        .I1(alu_io_in2[51]),
        .I2(ex_ctrl_alu_fn),
        .O(core__455_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2552" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__456
       (.I0(alu_io_in1[54]),
        .I1(alu_io_in2[54]),
        .I2(ex_ctrl_alu_fn),
        .O(core__456_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2543" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__457
       (.I0(alu_io_in1[57]),
        .I1(alu_io_in2[57]),
        .I2(ex_ctrl_alu_fn),
        .O(core__457_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2547" *) 
  LUT3 #(
    .INIT(8'h96)) 
    core__458
       (.I0(alu_io_in1[60]),
        .I1(alu_io_in2[60]),
        .I2(ex_ctrl_alu_fn),
        .O(core__458_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core__459
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core__459_n_0));
  LUT6 #(
    .INIT(64'hEE0E0000EE0EEE0E)) 
    core__46
       (.I0(core__56_n_0),
        .I1(frontend_n_386),
        .I2(frontend_n_404),
        .I3(frontend_n_393),
        .I4(frontend_n_395),
        .I5(frontend_n_409),
        .O(core__46_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2551" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    core__460
       (.I0(core_n_957),
        .I1(core_n_902),
        .I2(core__117_n_0),
        .O(core__460_n_0));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__461
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [39]),
        .I3(csr_io_tval),
        .O(\csr/p_1_in [39]));
  CARRY4 core__461_i_10
       (.CI(\<const0> ),
        .CO({core__461_i_10_n_0,core__461_i_10_n_1,core__461_i_10_n_2,core__461_i_10_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1697,core_n_1698,core_n_1699,core_n_1700}));
  CARRY4 core__461_i_3
       (.CI(core__461_i_5_n_0),
        .CO(_T_2520),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,core_n_1696}));
  CARRY4 core__461_i_4
       (.CI(core__461_i_7_n_0),
        .CO(_T_2522),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,core_n_652}));
  CARRY4 core__461_i_5
       (.CI(core__461_i_9_n_0),
        .CO({core__461_i_5_n_0,core__461_i_5_n_1,core__461_i_5_n_2,core__461_i_5_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core__315_n_0,core__314_n_0,core__313_n_0,core__312_n_0}));
  CARRY4 core__461_i_7
       (.CI(core__461_i_10_n_0),
        .CO({core__461_i_7_n_0,core__461_i_7_n_1,core__461_i_7_n_2,core__461_i_7_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1701,core_n_1702,core_n_1703,core_n_1704}));
  CARRY4 core__461_i_9
       (.CI(\<const0> ),
        .CO({core__461_i_9_n_0,core__461_i_9_n_1,core__461_i_9_n_2,core__461_i_9_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core__311_n_0,core__310_n_0,core__309_n_0,core__308_n_0}));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__462
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [30]),
        .I3(core_n_976),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [30]));
  CARRY4 core__462_i_10
       (.CI(\<const0> ),
        .CO({_T_2431,core__462_i_10_n_2,core__462_i_10_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,core_n_1795,core_n_1796,core_rep__36_n_0}));
  CARRY4 core__462_i_11
       (.CI(\<const0> ),
        .CO({_T_2428,core__462_i_11_n_2,core__462_i_11_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,core_n_1793,core_n_1794,core_rep__35_n_0}));
  CARRY4 core__462_i_12
       (.CI(\<const0> ),
        .CO({_T_2498,core__462_i_12_n_2,core__462_i_12_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,core_n_1788,core_n_1789,core__198_n_0}));
  CARRY4 core__462_i_3
       (.CI(\<const0> ),
        .CO({_T_2437,core__462_i_3_n_2,core__462_i_3_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,core_n_1797,core_n_1798,core__199_n_0}));
  CARRY4 core__462_i_4
       (.CI(\<const0> ),
        .CO({_T_2504,core__462_i_4_n_2,core__462_i_4_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,core_n_1338,core_n_1339,core_n_1340}));
  CARRY4 core__462_i_5
       (.CI(\<const0> ),
        .CO({_T_2507,core__462_i_5_n_2,core__462_i_5_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,core_n_1790,core_n_1791,core_n_1792}));
  CARRY4 core__462_i_6
       (.CI(\<const0> ),
        .CO({_T_2422,core__462_i_6_n_2,core__462_i_6_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,core_n_1332,core_n_1333,core_n_1334}));
  CARRY4 core__462_i_7
       (.CI(\<const0> ),
        .CO({_T_2499,core__462_i_7_n_2,core__462_i_7_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,core_n_1335,core_n_1336,core_n_1337}));
  CARRY4 core__462_i_8
       (.CI(\<const0> ),
        .CO({_T_2434,core__462_i_8_n_2,core__462_i_8_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,core_n_1341,core_n_1342,core__197_n_0}));
  CARRY4 core__462_i_9
       (.CI(\<const0> ),
        .CO({_T_2425,core__462_i_9_n_2,core__462_i_9_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,core_n_1783,core_n_1784,core_n_1785}));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__463
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [31]),
        .I3(core_n_975),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [31]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__464
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [32]),
        .I3(core_n_974),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [32]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__465
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [33]),
        .I3(core_n_973),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [33]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__466
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [34]),
        .I3(core_n_972),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [34]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__467
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [35]),
        .I3(core_n_971),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [35]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__468
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [36]),
        .I3(core_n_970),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [36]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__469
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [37]),
        .I3(core_n_969),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [37]));
  LUT6 #(
    .INIT(64'h0000010000001111)) 
    core__47
       (.I0(frontend_n_389),
        .I1(_T_1050[2]),
        .I2(_T_1005[4]),
        .I3(_T_1031[14]),
        .I4(_T_1031[3]),
        .I5(frontend_n_396),
        .O(core__47_n_0));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__470
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [38]),
        .I3(core_n_968),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [38]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__471
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [5]),
        .I3(core_n_966),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [5]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__472
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_5044 [4]),
        .I3(core_n_965),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [4]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__473
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_5044 [3]),
        .I3(core_n_964),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [3]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__474
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_5044 [2]),
        .I3(core_n_962),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [2]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__475
       (.I0(core_n_957),
        .I1(core_n_902),
        .I2(\csr/_T_5044 [1]),
        .I3(core_n_959),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [1]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__476
       (.I0(core_n_957),
        .I1(core_n_902),
        .I2(\csr/_T_5044 [0]),
        .I3(core_n_958),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [0]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__477
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [29]),
        .I3(core_n_956),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [29]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__478
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [28]),
        .I3(core_n_955),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [28]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__479
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [27]),
        .I3(core_n_954),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [27]));
  LUT6 #(
    .INIT(64'h41000041FFFFFFFF)) 
    core__48
       (.I0(dcache_n_551),
        .I1(dcache_n_550),
        .I2(ibuf_io_inst_0_bits_inst_rd[2]),
        .I3(dcache_n_542),
        .I4(ibuf_io_inst_0_bits_inst_rd[3]),
        .I5(frontend_n_376),
        .O(core__48_n_0));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__480
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [26]),
        .I3(core_n_953),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [26]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__481
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [25]),
        .I3(core_n_952),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [25]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__482
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [24]),
        .I3(core_n_951),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [24]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__483
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [23]),
        .I3(core_n_950),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [23]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__484
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [22]),
        .I3(core_n_949),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [22]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__485
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [21]),
        .I3(core_n_948),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [21]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__486
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [20]),
        .I3(core_n_946),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [20]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__487
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [19]),
        .I3(core_n_945),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [19]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__488
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [18]),
        .I3(core_n_944),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [18]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__489
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [17]),
        .I3(core_n_943),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [17]));
  LUT2 #(
    .INIT(4'h1)) 
    core__49
       (.I0(frontend_n_232),
        .I1(core_n_1102),
        .O(core__49_n_0));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__490
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [16]),
        .I3(core_n_942),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [16]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__491
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [15]),
        .I3(core_n_941),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [15]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__492
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [14]),
        .I3(core_n_940),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [14]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__493
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [13]),
        .I3(core_n_914),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [13]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__494
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [11]),
        .I3(core_n_913),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [11]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__495
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [10]),
        .I3(core_n_912),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [10]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__496
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [9]),
        .I3(core_n_910),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [9]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__497
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [8]),
        .I3(core_n_908),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [8]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__498
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [6]),
        .I3(core_n_906),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [6]));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__499
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [7]),
        .I3(core_n_904),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [7]));
  LUT6 #(
    .INIT(64'h3FAA33AA3FAA3FAA)) 
    core__5
       (.I0(core_n_16),
        .I1(frontend_n_265),
        .I2(frontend_n_419),
        .I3(_T_1790),
        .I4(core_n_1256),
        .I5(frontend_n_352),
        .O(core__5_n_0));
  LUT6 #(
    .INIT(64'h5555555555555554)) 
    core__50
       (.I0(ibuf_io_inst_0_bits_raw[12]),
        .I1(ibuf_io_inst_0_bits_raw[3]),
        .I2(ibuf_io_inst_0_bits_raw[4]),
        .I3(ibuf_io_inst_0_bits_raw[2]),
        .I4(ibuf_io_inst_0_bits_raw[5]),
        .I5(ibuf_io_inst_0_bits_raw[6]),
        .O(core__50_n_0));
  LUT5 #(
    .INIT(32'h2020FD20)) 
    core__500
       (.I0(core_n_1020),
        .I1(core_n_902),
        .I2(\csr/_T_4899 [12]),
        .I3(core_n_897),
        .I4(dcache_n_558),
        .O(\csr/p_1_in [12]));
  LUT6 #(
    .INIT(64'h5511151544000404)) 
    core__501
       (.I0(target_reset),
        .I1(\csr/reg_mstatus_mie ),
        .I2(core_n_1005),
        .I3(\csr/_T_4899 [7]),
        .I4(core_n_1008),
        .I5(core_n_86),
        .O(core__501_n_0));
  LUT6 #(
    .INIT(64'hFBFBFFBBEAEAEEAA)) 
    core__502
       (.I0(target_reset),
        .I1(\csr/reg_mstatus_mie ),
        .I2(\csr/_T_4899 [11]),
        .I3(core_n_1007),
        .I4(core_n_1008),
        .I5(core_n_1002),
        .O(core__502_n_0));
  LUT6 #(
    .INIT(64'hFBFBFFBBEAEAEEAA)) 
    core__503
       (.I0(target_reset),
        .I1(\csr/reg_mstatus_mie ),
        .I2(\csr/_T_4899 [12]),
        .I3(core_n_1006),
        .I4(core_n_1008),
        .I5(core_n_901),
        .O(core__503_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2501" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    core__504
       (.I0(core_n_1020),
        .I1(core_n_963),
        .I2(core__117_n_0),
        .O(core__504_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2501" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__505
       (.I0(core_n_1020),
        .I1(core_n_963),
        .I2(\csr/_T_5044 [63]),
        .I3(core_n_1014),
        .O(core__505_n_0));
  LUT4 #(
    .INIT(16'h20FD)) 
    core__506
       (.I0(core_n_1020),
        .I1(core_n_963),
        .I2(\csr/_T_5044 [3]),
        .I3(core_n_1012),
        .O(core__506_n_0));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__507
       (.I0(core_n_1020),
        .I1(core_n_963),
        .I2(\csr/_T_5044 [2]),
        .I3(core__433_n_0),
        .O(core__507_n_0));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__508
       (.I0(core_n_1020),
        .I1(core_n_963),
        .I2(\csr/_T_5044 [1]),
        .I3(core_n_1016),
        .O(core__508_n_0));
  LUT4 #(
    .INIT(16'h20FD)) 
    core__509
       (.I0(core_n_1020),
        .I1(core_n_963),
        .I2(\csr/_T_5044 [0]),
        .I3(core__119_n_0),
        .O(core__509_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    core__51
       (.I0(frontend_n_404),
        .I1(_T_1005[4]),
        .O(core__51_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2503" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    core__510
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(core__117_n_0),
        .O(core__510_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2491" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__511
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [39]),
        .I3(wb_reg_pc[39]),
        .O(\csr/_GEN_350 [39]));
  (* SOFT_HLUTNM = "soft_lutpair2515" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__512
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [30]),
        .I3(wb_reg_pc[30]),
        .O(\csr/_GEN_350 [30]));
  (* SOFT_HLUTNM = "soft_lutpair2506" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__513
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [31]),
        .I3(wb_reg_pc[31]),
        .O(\csr/_GEN_350 [31]));
  (* SOFT_HLUTNM = "soft_lutpair2513" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__514
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [32]),
        .I3(wb_reg_pc[32]),
        .O(\csr/_GEN_350 [32]));
  (* SOFT_HLUTNM = "soft_lutpair2510" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__515
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [33]),
        .I3(wb_reg_pc[33]),
        .O(\csr/_GEN_350 [33]));
  (* SOFT_HLUTNM = "soft_lutpair2526" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__516
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [34]),
        .I3(wb_reg_pc[34]),
        .O(\csr/_GEN_350 [34]));
  (* SOFT_HLUTNM = "soft_lutpair2531" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__517
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [35]),
        .I3(wb_reg_pc[35]),
        .O(\csr/_GEN_350 [35]));
  (* SOFT_HLUTNM = "soft_lutpair2514" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__518
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [36]),
        .I3(wb_reg_pc[36]),
        .O(\csr/_GEN_350 [36]));
  (* SOFT_HLUTNM = "soft_lutpair2532" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__519
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [37]),
        .I3(wb_reg_pc[37]),
        .O(\csr/_GEN_350 [37]));
  (* SOFT_HLUTNM = "soft_lutpair2485" *) 
  LUT5 #(
    .INIT(32'hFFFFFF08)) 
    core__52
       (.I0(ibuf_io_inst_0_bits_raw[12]),
        .I1(frontend_n_294),
        .I2(frontend_n_293),
        .I3(frontend_n_285),
        .I4(ibuf_io_inst_0_bits_raw[1]),
        .O(core__52_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2504" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__520
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [38]),
        .I3(wb_reg_pc[38]),
        .O(\csr/_GEN_350 [38]));
  (* SOFT_HLUTNM = "soft_lutpair2503" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__521
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [5]),
        .I3(wb_reg_pc[5]),
        .O(\csr/_GEN_350 [5]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__522
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_5044 [4]),
        .I3(wb_reg_pc[4]),
        .O(\csr/_GEN_350 [4]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__523
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_5044 [3]),
        .I3(wb_reg_pc[3]),
        .O(\csr/_GEN_350 [3]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__524
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_5044 [2]),
        .I3(wb_reg_pc[2]),
        .O(\csr/_GEN_350 [2]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__525
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_5044 [1]),
        .I3(wb_reg_pc[1]),
        .O(\csr/_GEN_350 [1]));
  (* SOFT_HLUTNM = "soft_lutpair2533" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__526
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [29]),
        .I3(wb_reg_pc[29]),
        .O(\csr/_GEN_350 [29]));
  (* SOFT_HLUTNM = "soft_lutpair2534" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__527
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [28]),
        .I3(wb_reg_pc[28]),
        .O(\csr/_GEN_350 [28]));
  (* SOFT_HLUTNM = "soft_lutpair2511" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__528
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [27]),
        .I3(wb_reg_pc[27]),
        .O(\csr/_GEN_350 [27]));
  (* SOFT_HLUTNM = "soft_lutpair2512" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__529
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [26]),
        .I3(wb_reg_pc[26]),
        .O(\csr/_GEN_350 [26]));
  (* SOFT_HLUTNM = "soft_lutpair2485" *) 
  LUT3 #(
    .INIT(8'h40)) 
    core__53
       (.I0(frontend_n_293),
        .I1(frontend_n_294),
        .I2(ibuf_io_inst_0_bits_raw[12]),
        .O(core__53_n_0));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__530
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [25]),
        .I3(wb_reg_pc[25]),
        .O(\csr/_GEN_350 [25]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__531
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [24]),
        .I3(wb_reg_pc[24]),
        .O(\csr/_GEN_350 [24]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__532
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [23]),
        .I3(wb_reg_pc[23]),
        .O(\csr/_GEN_350 [23]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__533
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [22]),
        .I3(wb_reg_pc[22]),
        .O(\csr/_GEN_350 [22]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__534
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [21]),
        .I3(wb_reg_pc[21]),
        .O(\csr/_GEN_350 [21]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__535
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [20]),
        .I3(wb_reg_pc[20]),
        .O(\csr/_GEN_350 [20]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__536
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [19]),
        .I3(wb_reg_pc[19]),
        .O(\csr/_GEN_350 [19]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__537
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [18]),
        .I3(wb_reg_pc[18]),
        .O(\csr/_GEN_350 [18]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__538
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [17]),
        .I3(wb_reg_pc[17]),
        .O(\csr/_GEN_350 [17]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__539
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [16]),
        .I3(wb_reg_pc[16]),
        .O(\csr/_GEN_350 [16]));
  LUT6 #(
    .INIT(64'h5555555515555555)) 
    core__54
       (.I0(ibuf_io_inst_0_bits_raw[2]),
        .I1(frontend_n_304),
        .I2(ibuf_io_inst_0_bits_raw[12]),
        .I3(frontend_n_269),
        .I4(core__80_n_0),
        .I5(ibuf_io_inst_0_bits_raw[14]),
        .O(core__54_n_0));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__540
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [15]),
        .I3(wb_reg_pc[15]),
        .O(\csr/_GEN_350 [15]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__541
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [14]),
        .I3(wb_reg_pc[14]),
        .O(\csr/_GEN_350 [14]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__542
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [13]),
        .I3(wb_reg_pc[13]),
        .O(\csr/_GEN_350 [13]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__543
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [11]),
        .I3(wb_reg_pc[11]),
        .O(\csr/_GEN_350 [11]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__544
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [10]),
        .I3(wb_reg_pc[10]),
        .O(\csr/_GEN_350 [10]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__545
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [9]),
        .I3(wb_reg_pc[9]),
        .O(\csr/_GEN_350 [9]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__546
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [8]),
        .I3(wb_reg_pc[8]),
        .O(\csr/_GEN_350 [8]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__547
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [6]),
        .I3(wb_reg_pc[6]),
        .O(\csr/_GEN_350 [6]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__548
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [7]),
        .I3(wb_reg_pc[7]),
        .O(\csr/_GEN_350 [7]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__549
       (.I0(core_n_1020),
        .I1(core_n_909),
        .I2(\csr/_T_4899 [12]),
        .I3(wb_reg_pc[12]),
        .O(\csr/_GEN_350 [12]));
  (* SOFT_HLUTNM = "soft_lutpair2545" *) 
  LUT3 #(
    .INIT(8'h10)) 
    core__55
       (.I0(_T_1005[4]),
        .I1(_T_1031[3]),
        .I2(_T_1050[2]),
        .O(core__55_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2551" *) 
  LUT3 #(
    .INIT(8'h20)) 
    core__550
       (.I0(core_n_957),
        .I1(core__113_n_0),
        .I2(\csr/_T_5044 [0]),
        .O(core__550_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2502" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    core__551
       (.I0(core_n_895),
        .I1(core_n_995),
        .I2(core_n_992),
        .O(core__551_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2502" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__552
       (.I0(core_n_895),
        .I1(core_n_995),
        .I2(\csr/_T_5044 [63]),
        .I3(core_n_1014),
        .O(core__552_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2505" *) 
  LUT3 #(
    .INIT(8'h20)) 
    core__553
       (.I0(core_n_895),
        .I1(core_n_995),
        .I2(\csr/_T_5044 [4]),
        .O(core__553_n_0));
  LUT4 #(
    .INIT(16'h20FD)) 
    core__554
       (.I0(core_n_895),
        .I1(core_n_995),
        .I2(\csr/_T_5044 [3]),
        .I3(core_n_1012),
        .O(core__554_n_0));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__555
       (.I0(core_n_895),
        .I1(core_n_995),
        .I2(\csr/_T_5044 [2]),
        .I3(core__433_n_0),
        .O(core__555_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2505" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__556
       (.I0(core_n_895),
        .I1(core_n_995),
        .I2(\csr/_T_5044 [1]),
        .I3(core_n_1016),
        .O(core__556_n_0));
  LUT4 #(
    .INIT(16'h20FD)) 
    core__557
       (.I0(core_n_895),
        .I1(core_n_995),
        .I2(\csr/_T_5044 [0]),
        .I3(core__119_n_0),
        .O(core__557_n_0));
  LUT3 #(
    .INIT(8'hF2)) 
    core__558
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(core_n_992),
        .O(core__558_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2491" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__559
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [39]),
        .I3(wb_reg_pc[39]),
        .O(\csr/_GEN_369 [39]));
  (* SOFT_HLUTNM = "soft_lutpair2545" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    core__56
       (.I0(_T_1005[4]),
        .I1(_T_1050[2]),
        .I2(_T_1050[5]),
        .O(core__56_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2515" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__560
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [30]),
        .I3(wb_reg_pc[30]),
        .O(\csr/_GEN_369 [30]));
  (* SOFT_HLUTNM = "soft_lutpair2506" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__561
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [31]),
        .I3(wb_reg_pc[31]),
        .O(\csr/_GEN_369 [31]));
  (* SOFT_HLUTNM = "soft_lutpair2513" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__562
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [32]),
        .I3(wb_reg_pc[32]),
        .O(\csr/_GEN_369 [32]));
  (* SOFT_HLUTNM = "soft_lutpair2510" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__563
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [33]),
        .I3(wb_reg_pc[33]),
        .O(\csr/_GEN_369 [33]));
  (* SOFT_HLUTNM = "soft_lutpair2526" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__564
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [34]),
        .I3(wb_reg_pc[34]),
        .O(\csr/_GEN_369 [34]));
  (* SOFT_HLUTNM = "soft_lutpair2531" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__565
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [35]),
        .I3(wb_reg_pc[35]),
        .O(\csr/_GEN_369 [35]));
  (* SOFT_HLUTNM = "soft_lutpair2514" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__566
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [36]),
        .I3(wb_reg_pc[36]),
        .O(\csr/_GEN_369 [36]));
  (* SOFT_HLUTNM = "soft_lutpair2532" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__567
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [37]),
        .I3(wb_reg_pc[37]),
        .O(\csr/_GEN_369 [37]));
  (* SOFT_HLUTNM = "soft_lutpair2504" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__568
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [38]),
        .I3(wb_reg_pc[38]),
        .O(\csr/_GEN_369 [38]));
  (* SOFT_HLUTNM = "soft_lutpair2516" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__569
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [5]),
        .I3(wb_reg_pc[5]),
        .O(\csr/_GEN_369 [5]));
  LUT6 #(
    .INIT(64'hFDDD0000FFFFFFFF)) 
    core__57
       (.I0(core__80_n_0),
        .I1(ibuf_io_inst_0_bits_raw[14]),
        .I2(ibuf_io_inst_0_bits_raw[12]),
        .I3(frontend_n_304),
        .I4(frontend_n_312),
        .I5(frontend_n_300),
        .O(core__57_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2541" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__570
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_5044 [4]),
        .I3(wb_reg_pc[4]),
        .O(\csr/_GEN_369 [4]));
  (* SOFT_HLUTNM = "soft_lutpair2517" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__571
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_5044 [3]),
        .I3(wb_reg_pc[3]),
        .O(\csr/_GEN_369 [3]));
  (* SOFT_HLUTNM = "soft_lutpair2507" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__572
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_5044 [2]),
        .I3(wb_reg_pc[2]),
        .O(\csr/_GEN_369 [2]));
  (* SOFT_HLUTNM = "soft_lutpair2518" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__573
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_5044 [1]),
        .I3(wb_reg_pc[1]),
        .O(\csr/_GEN_369 [1]));
  (* SOFT_HLUTNM = "soft_lutpair2533" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__574
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [29]),
        .I3(wb_reg_pc[29]),
        .O(\csr/_GEN_369 [29]));
  (* SOFT_HLUTNM = "soft_lutpair2534" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__575
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [28]),
        .I3(wb_reg_pc[28]),
        .O(\csr/_GEN_369 [28]));
  (* SOFT_HLUTNM = "soft_lutpair2511" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__576
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [27]),
        .I3(wb_reg_pc[27]),
        .O(\csr/_GEN_369 [27]));
  (* SOFT_HLUTNM = "soft_lutpair2512" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__577
       (.I0(core_n_1020),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [26]),
        .I3(wb_reg_pc[26]),
        .O(\csr/_GEN_369 [26]));
  (* SOFT_HLUTNM = "soft_lutpair2524" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__578
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [25]),
        .I3(wb_reg_pc[25]),
        .O(\csr/_GEN_369 [25]));
  (* SOFT_HLUTNM = "soft_lutpair2525" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__579
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [24]),
        .I3(wb_reg_pc[24]),
        .O(\csr/_GEN_369 [24]));
  LUT6 #(
    .INIT(64'h04000000FFFFFFFF)) 
    core__58
       (.I0(ibuf_io_inst_0_bits_raw[12]),
        .I1(core__80_n_0),
        .I2(core__73_n_0),
        .I3(ibuf_io_inst_0_bits_raw[15]),
        .I4(frontend_n_304),
        .I5(frontend_n_300),
        .O(core__58_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2536" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__580
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [23]),
        .I3(wb_reg_pc[23]),
        .O(\csr/_GEN_369 [23]));
  (* SOFT_HLUTNM = "soft_lutpair2519" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__581
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [22]),
        .I3(wb_reg_pc[22]),
        .O(\csr/_GEN_369 [22]));
  (* SOFT_HLUTNM = "soft_lutpair2537" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__582
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [21]),
        .I3(wb_reg_pc[21]),
        .O(\csr/_GEN_369 [21]));
  (* SOFT_HLUTNM = "soft_lutpair2538" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__583
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [20]),
        .I3(wb_reg_pc[20]),
        .O(\csr/_GEN_369 [20]));
  (* SOFT_HLUTNM = "soft_lutpair2542" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__584
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [19]),
        .I3(wb_reg_pc[19]),
        .O(\csr/_GEN_369 [19]));
  (* SOFT_HLUTNM = "soft_lutpair2539" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__585
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [18]),
        .I3(wb_reg_pc[18]),
        .O(\csr/_GEN_369 [18]));
  (* SOFT_HLUTNM = "soft_lutpair2520" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__586
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [17]),
        .I3(wb_reg_pc[17]),
        .O(\csr/_GEN_369 [17]));
  (* SOFT_HLUTNM = "soft_lutpair2540" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__587
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [16]),
        .I3(wb_reg_pc[16]),
        .O(\csr/_GEN_369 [16]));
  (* SOFT_HLUTNM = "soft_lutpair2521" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__588
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [15]),
        .I3(wb_reg_pc[15]),
        .O(\csr/_GEN_369 [15]));
  (* SOFT_HLUTNM = "soft_lutpair2530" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__589
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [14]),
        .I3(wb_reg_pc[14]),
        .O(\csr/_GEN_369 [14]));
  LUT6 #(
    .INIT(64'h0400000000000000)) 
    core__59
       (.I0(ibuf_io_inst_0_bits_raw[12]),
        .I1(core__80_n_0),
        .I2(core__73_n_0),
        .I3(ibuf_io_inst_0_bits_raw[15]),
        .I4(frontend_n_304),
        .I5(frontend_n_300),
        .O(core__59_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2522" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__590
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [13]),
        .I3(wb_reg_pc[13]),
        .O(\csr/_GEN_369 [13]));
  (* SOFT_HLUTNM = "soft_lutpair2529" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__591
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [11]),
        .I3(wb_reg_pc[11]),
        .O(\csr/_GEN_369 [11]));
  (* SOFT_HLUTNM = "soft_lutpair2508" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__592
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [10]),
        .I3(wb_reg_pc[10]),
        .O(\csr/_GEN_369 [10]));
  (* SOFT_HLUTNM = "soft_lutpair2523" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__593
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [9]),
        .I3(wb_reg_pc[9]),
        .O(\csr/_GEN_369 [9]));
  (* SOFT_HLUTNM = "soft_lutpair2528" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__594
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [8]),
        .I3(wb_reg_pc[8]),
        .O(\csr/_GEN_369 [8]));
  (* SOFT_HLUTNM = "soft_lutpair2527" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__595
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [6]),
        .I3(wb_reg_pc[6]),
        .O(\csr/_GEN_369 [6]));
  (* SOFT_HLUTNM = "soft_lutpair2509" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__596
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [7]),
        .I3(wb_reg_pc[7]),
        .O(\csr/_GEN_369 [7]));
  (* SOFT_HLUTNM = "soft_lutpair2535" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__597
       (.I0(core_n_895),
        .I1(core_n_907),
        .I2(\csr/_T_4899 [12]),
        .I3(wb_reg_pc[12]),
        .O(\csr/_GEN_369 [12]));
  (* SOFT_HLUTNM = "soft_lutpair2492" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    core__598
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/reg_dcsr_prv ),
        .O(core__598_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2492" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__599
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [39]),
        .I3(wb_reg_pc[39]),
        .O(\csr/_GEN_364 [39]));
  LUT6 #(
    .INIT(64'hFFFFCFFFAAAAAAAA)) 
    core__6
       (.I0(core_n_0),
        .I1(id_ctrl_alu_dw),
        .I2(frontend_n_352),
        .I3(frontend_n_355),
        .I4(core_n_1089),
        .I5(_T_1790),
        .O(core__6_n_0));
  LUT5 #(
    .INIT(32'h20000000)) 
    core__60
       (.I0(frontend_n_269),
        .I1(ibuf_io_inst_0_bits_raw[14]),
        .I2(frontend_n_268),
        .I3(ibuf_io_inst_0_bits_raw[11]),
        .I4(ibuf_io_inst_0_bits_raw[12]),
        .O(core__60_n_0));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__600
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [30]),
        .I3(wb_reg_pc[30]),
        .O(\csr/_GEN_364 [30]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__601
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [31]),
        .I3(wb_reg_pc[31]),
        .O(\csr/_GEN_364 [31]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__602
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [32]),
        .I3(wb_reg_pc[32]),
        .O(\csr/_GEN_364 [32]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__603
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [33]),
        .I3(wb_reg_pc[33]),
        .O(\csr/_GEN_364 [33]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__604
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [34]),
        .I3(wb_reg_pc[34]),
        .O(\csr/_GEN_364 [34]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__605
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [35]),
        .I3(wb_reg_pc[35]),
        .O(\csr/_GEN_364 [35]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__606
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [36]),
        .I3(wb_reg_pc[36]),
        .O(\csr/_GEN_364 [36]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__607
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [37]),
        .I3(wb_reg_pc[37]),
        .O(\csr/_GEN_364 [37]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__608
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [38]),
        .I3(wb_reg_pc[38]),
        .O(\csr/_GEN_364 [38]));
  (* SOFT_HLUTNM = "soft_lutpair2516" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__609
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [5]),
        .I3(wb_reg_pc[5]),
        .O(\csr/_GEN_364 [5]));
  LUT6 #(
    .INIT(64'h1000100055551000)) 
    core__61
       (.I0(ibuf_io_inst_0_bits_raw[1]),
        .I1(core__67_n_0),
        .I2(ibuf_io_inst_0_bits_raw[0]),
        .I3(ibuf_io_inst_0_bits_raw[15]),
        .I4(frontend_n_285),
        .I5(ibuf_io_inst_0_bits_raw[12]),
        .O(core__61_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2541" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__610
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_5044 [4]),
        .I3(wb_reg_pc[4]),
        .O(\csr/_GEN_364 [4]));
  (* SOFT_HLUTNM = "soft_lutpair2517" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__611
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_5044 [3]),
        .I3(wb_reg_pc[3]),
        .O(\csr/_GEN_364 [3]));
  (* SOFT_HLUTNM = "soft_lutpair2507" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__612
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_5044 [2]),
        .I3(wb_reg_pc[2]),
        .O(\csr/_GEN_364 [2]));
  (* SOFT_HLUTNM = "soft_lutpair2518" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__613
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_5044 [1]),
        .I3(wb_reg_pc[1]),
        .O(\csr/_GEN_364 [1]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__614
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [29]),
        .I3(wb_reg_pc[29]),
        .O(\csr/_GEN_364 [29]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__615
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [28]),
        .I3(wb_reg_pc[28]),
        .O(\csr/_GEN_364 [28]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__616
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [27]),
        .I3(wb_reg_pc[27]),
        .O(\csr/_GEN_364 [27]));
  LUT4 #(
    .INIT(16'hFD20)) 
    core__617
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [26]),
        .I3(wb_reg_pc[26]),
        .O(\csr/_GEN_364 [26]));
  (* SOFT_HLUTNM = "soft_lutpair2524" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__618
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [25]),
        .I3(wb_reg_pc[25]),
        .O(\csr/_GEN_364 [25]));
  (* SOFT_HLUTNM = "soft_lutpair2525" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__619
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [24]),
        .I3(wb_reg_pc[24]),
        .O(\csr/_GEN_364 [24]));
  LUT6 #(
    .INIT(64'h00ACFFAC00A000A0)) 
    core__62
       (.I0(ibuf_io_inst_0_bits_raw[3]),
        .I1(core__77_n_0),
        .I2(frontend_n_267),
        .I3(ibuf_io_inst_0_bits_raw[1]),
        .I4(frontend_n_318),
        .I5(ibuf_io_inst_0_bits_raw[8]),
        .O(core__62_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2536" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__620
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [23]),
        .I3(wb_reg_pc[23]),
        .O(\csr/_GEN_364 [23]));
  (* SOFT_HLUTNM = "soft_lutpair2519" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__621
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [22]),
        .I3(wb_reg_pc[22]),
        .O(\csr/_GEN_364 [22]));
  (* SOFT_HLUTNM = "soft_lutpair2537" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__622
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [21]),
        .I3(wb_reg_pc[21]),
        .O(\csr/_GEN_364 [21]));
  (* SOFT_HLUTNM = "soft_lutpair2538" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__623
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [20]),
        .I3(wb_reg_pc[20]),
        .O(\csr/_GEN_364 [20]));
  (* SOFT_HLUTNM = "soft_lutpair2542" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__624
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [19]),
        .I3(wb_reg_pc[19]),
        .O(\csr/_GEN_364 [19]));
  (* SOFT_HLUTNM = "soft_lutpair2539" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__625
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [18]),
        .I3(wb_reg_pc[18]),
        .O(\csr/_GEN_364 [18]));
  (* SOFT_HLUTNM = "soft_lutpair2520" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__626
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [17]),
        .I3(wb_reg_pc[17]),
        .O(\csr/_GEN_364 [17]));
  (* SOFT_HLUTNM = "soft_lutpair2540" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__627
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [16]),
        .I3(wb_reg_pc[16]),
        .O(\csr/_GEN_364 [16]));
  (* SOFT_HLUTNM = "soft_lutpair2521" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__628
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [15]),
        .I3(wb_reg_pc[15]),
        .O(\csr/_GEN_364 [15]));
  (* SOFT_HLUTNM = "soft_lutpair2530" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__629
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [14]),
        .I3(wb_reg_pc[14]),
        .O(\csr/_GEN_364 [14]));
  LUT6 #(
    .INIT(64'h00000200FFFFFFFF)) 
    core__63
       (.I0(ibuf_io_inst_0_bits_raw[9]),
        .I1(ibuf_io_inst_0_bits_raw[15]),
        .I2(ibuf_io_inst_0_bits_raw[14]),
        .I3(frontend_n_269),
        .I4(ibuf_io_inst_0_bits_raw[0]),
        .I5(ibuf_io_inst_0_bits_raw[1]),
        .O(core__63_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2522" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__630
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [13]),
        .I3(wb_reg_pc[13]),
        .O(\csr/_GEN_364 [13]));
  (* SOFT_HLUTNM = "soft_lutpair2529" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__631
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [11]),
        .I3(wb_reg_pc[11]),
        .O(\csr/_GEN_364 [11]));
  (* SOFT_HLUTNM = "soft_lutpair2508" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__632
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [10]),
        .I3(wb_reg_pc[10]),
        .O(\csr/_GEN_364 [10]));
  (* SOFT_HLUTNM = "soft_lutpair2523" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__633
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [9]),
        .I3(wb_reg_pc[9]),
        .O(\csr/_GEN_364 [9]));
  (* SOFT_HLUTNM = "soft_lutpair2528" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__634
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [8]),
        .I3(wb_reg_pc[8]),
        .O(\csr/_GEN_364 [8]));
  (* SOFT_HLUTNM = "soft_lutpair2527" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__635
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [6]),
        .I3(wb_reg_pc[6]),
        .O(\csr/_GEN_364 [6]));
  (* SOFT_HLUTNM = "soft_lutpair2509" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__636
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [7]),
        .I3(wb_reg_pc[7]),
        .O(\csr/_GEN_364 [7]));
  (* SOFT_HLUTNM = "soft_lutpair2535" *) 
  LUT4 #(
    .INIT(16'hFD20)) 
    core__637
       (.I0(core_n_895),
        .I1(core_n_947),
        .I2(\csr/_T_4899 [12]),
        .I3(wb_reg_pc[12]),
        .O(\csr/_GEN_364 [12]));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    core__638
       (.I0(core_n_2286),
        .I1(alu_io_in2[1]),
        .I2(core_n_2281),
        .I3(alu_io_in2[0]),
        .I4(core_n_2283),
        .I5(core__644_n_0),
        .O(core__638_n_0));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    core__639
       (.I0(core_n_2287),
        .I1(alu_io_in2[3]),
        .I2(core_n_2264),
        .I3(alu_io_in2[2]),
        .I4(core_n_2272),
        .I5(core_n_2255),
        .O(core__639_n_0));
  LUT6 #(
    .INIT(64'h00ACFFAC00A000A0)) 
    core__64
       (.I0(ibuf_io_inst_0_bits_raw[4]),
        .I1(core__77_n_0),
        .I2(frontend_n_267),
        .I3(ibuf_io_inst_0_bits_raw[1]),
        .I4(frontend_n_318),
        .I5(ibuf_io_inst_0_bits_raw[9]),
        .O(core__64_n_0));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    core__640
       (.I0(\alu/shin [63]),
        .I1(\alu/shamt ),
        .I2(\alu/shin [31]),
        .I3(alu_io_in2[4]),
        .I4(\alu/shin [47]),
        .I5(\alu/shin [15]),
        .O(core__640_n_0));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    core__641
       (.I0(core_n_2290),
        .I1(alu_io_in2[3]),
        .I2(core_n_2266),
        .I3(alu_io_in2[2]),
        .I4(core_n_2274),
        .I5(core_n_2257),
        .O(core__641_n_0));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    core__642
       (.I0(core_n_2288),
        .I1(alu_io_in2[1]),
        .I2(core_n_2286),
        .I3(core__645_n_0),
        .I4(core_n_2285),
        .I5(alu_io_in2[0]),
        .O(core__642_n_0));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    core__643
       (.I0(core_n_2292),
        .I1(alu_io_in2[3]),
        .I2(core_n_2268),
        .I3(alu_io_in2[2]),
        .I4(core_n_2276),
        .I5(core_n_2260),
        .O(core__643_n_0));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    core__644
       (.I0(core_n_2294),
        .I1(alu_io_in2[3]),
        .I2(core_n_2270),
        .I3(alu_io_in2[2]),
        .I4(core_n_2278),
        .I5(core_n_2262),
        .O(core__644_n_0));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    core__645
       (.I0(core_n_2289),
        .I1(alu_io_in2[3]),
        .I2(core_n_2274),
        .I3(core_n_2296),
        .I4(alu_io_in2[2]),
        .O(core__645_n_0));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    core__646
       (.I0(core_n_2291),
        .I1(alu_io_in2[3]),
        .I2(core_n_2276),
        .I3(core_n_2297),
        .I4(alu_io_in2[2]),
        .O(core__646_n_0));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    core__647
       (.I0(core_n_2293),
        .I1(alu_io_in2[3]),
        .I2(core_n_2278),
        .I3(core_n_2298),
        .I4(alu_io_in2[2]),
        .O(core__647_n_0));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    core__648
       (.I0(core_n_2295),
        .I1(alu_io_in2[3]),
        .I2(core_n_2287),
        .I3(core_n_2299),
        .I4(alu_io_in2[2]),
        .O(core__648_n_0));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    core__649
       (.I0(core_n_2303),
        .I1(alu_io_in2[1]),
        .I2(core_n_2301),
        .I3(alu_io_in2[0]),
        .I4(core_n_2302),
        .I5(core_n_2300),
        .O(core__649_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2479" *) 
  LUT5 #(
    .INIT(32'h15151555)) 
    core__65
       (.I0(ibuf_io_inst_0_bits_raw[1]),
        .I1(ibuf_io_inst_0_bits_raw[15]),
        .I2(ibuf_io_inst_0_bits_raw[0]),
        .I3(frontend_n_269),
        .I4(ibuf_io_inst_0_bits_raw[14]),
        .O(core__65_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__650
       (.I0(core_n_2304),
        .I1(alu_io_in2[1]),
        .I2(core_n_2302),
        .I3(core_n_2303),
        .I4(core_n_2301),
        .I5(alu_io_in2[0]),
        .O(core__650_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__651
       (.I0(core_n_2305),
        .I1(alu_io_in2[1]),
        .I2(core_n_2303),
        .I3(core_n_2304),
        .I4(core_n_2302),
        .I5(alu_io_in2[0]),
        .O(core__651_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__652
       (.I0(core_n_2306),
        .I1(alu_io_in2[1]),
        .I2(core_n_2304),
        .I3(core_n_2305),
        .I4(core_n_2303),
        .I5(alu_io_in2[0]),
        .O(core__652_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__653
       (.I0(core_n_2307),
        .I1(alu_io_in2[1]),
        .I2(core_n_2305),
        .I3(core_n_2306),
        .I4(core_n_2304),
        .I5(alu_io_in2[0]),
        .O(core__653_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__654
       (.I0(core_n_2308),
        .I1(alu_io_in2[1]),
        .I2(core_n_2306),
        .I3(core_n_2307),
        .I4(core_n_2305),
        .I5(alu_io_in2[0]),
        .O(core__654_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__655
       (.I0(core_n_2309),
        .I1(alu_io_in2[1]),
        .I2(core_n_2307),
        .I3(core_n_2308),
        .I4(core_n_2306),
        .I5(alu_io_in2[0]),
        .O(core__655_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__656
       (.I0(core_n_2310),
        .I1(alu_io_in2[1]),
        .I2(core_n_2308),
        .I3(core_n_2309),
        .I4(core_n_2307),
        .I5(alu_io_in2[0]),
        .O(core__656_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__657
       (.I0(core_n_2311),
        .I1(alu_io_in2[1]),
        .I2(core_n_2309),
        .I3(core_n_2310),
        .I4(core_n_2308),
        .I5(alu_io_in2[0]),
        .O(core__657_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__658
       (.I0(core_n_2312),
        .I1(alu_io_in2[1]),
        .I2(core_n_2310),
        .I3(core_n_2311),
        .I4(core_n_2309),
        .I5(alu_io_in2[0]),
        .O(core__658_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__659
       (.I0(core_n_2313),
        .I1(alu_io_in2[1]),
        .I2(core_n_2311),
        .I3(core_n_2312),
        .I4(core_n_2310),
        .I5(alu_io_in2[0]),
        .O(core__659_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2482" *) 
  LUT4 #(
    .INIT(16'hE000)) 
    core__66
       (.I0(ibuf_io_inst_0_bits_raw[14]),
        .I1(frontend_n_269),
        .I2(ibuf_io_inst_0_bits_raw[0]),
        .I3(ibuf_io_inst_0_bits_raw[15]),
        .O(core__66_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__660
       (.I0(core_n_2314),
        .I1(alu_io_in2[1]),
        .I2(core_n_2312),
        .I3(core_n_2313),
        .I4(core_n_2311),
        .I5(alu_io_in2[0]),
        .O(core__660_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__661
       (.I0(core_n_2316),
        .I1(alu_io_in2[1]),
        .I2(core_n_2313),
        .I3(core_n_2314),
        .I4(core_n_2312),
        .I5(alu_io_in2[0]),
        .O(core__661_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__662
       (.I0(core_n_2315),
        .I1(alu_io_in2[1]),
        .I2(core_n_2314),
        .I3(core_n_2316),
        .I4(core_n_2313),
        .I5(alu_io_in2[0]),
        .O(core__662_n_0));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    core__663
       (.I0(\alu/_T_121 ),
        .I1(alu_io_in2[1]),
        .I2(core_n_2316),
        .I3(core_n_2315),
        .I4(core_n_2314),
        .I5(alu_io_in2[0]),
        .O(core__663_n_0));
  LUT6 #(
    .INIT(64'h5454FE54FEFEFE54)) 
    core__664
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core__291_n_0),
        .I3(\div/_T_122 ),
        .I4(core__191_n_0),
        .I5(core_n_310),
        .O(core__664_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__665
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[23]),
        .I4(core_n_288),
        .O(core__665_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__666
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[22]),
        .I4(core_n_287),
        .O(core__666_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__667
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[21]),
        .I4(core_n_286),
        .O(core__667_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__668
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[19]),
        .I4(core_n_285),
        .O(core__668_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__669
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[18]),
        .I4(core_n_284),
        .O(core__669_n_0));
  LUT6 #(
    .INIT(64'h000000000407F4F7)) 
    core__67
       (.I0(frontend_io_cpu_resp_bits_data[30]),
        .I1(frontend_io_cpu_resp_bits_pc[1]),
        .I2(\ibuf/_T_100 ),
        .I3(frontend_io_cpu_resp_bits_data[14]),
        .I4(core_n_2087),
        .I5(frontend_n_269),
        .O(core__67_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__670
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[16]),
        .I4(core_n_283),
        .O(core__670_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__671
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[15]),
        .I4(core_n_282),
        .O(core__671_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__672
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[13]),
        .I4(core_n_281),
        .O(core__672_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__673
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[12]),
        .I4(core_n_280),
        .O(core__673_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__674
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[11]),
        .I4(core_n_279),
        .O(core__674_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__675
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[10]),
        .I4(core_n_278),
        .O(core__675_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__676
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[8]),
        .I4(core_n_277),
        .O(core__676_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__677
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[7]),
        .I4(core_n_276),
        .O(core__677_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__678
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[5]),
        .I4(core_n_275),
        .O(core__678_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__679
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[4]),
        .I4(core_n_274),
        .O(core__679_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2479" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    core__68
       (.I0(ibuf_io_inst_0_bits_raw[15]),
        .I1(ibuf_io_inst_0_bits_raw[14]),
        .I2(frontend_n_269),
        .I3(ibuf_io_inst_0_bits_raw[0]),
        .O(core__68_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__680
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[3]),
        .I4(core_n_273),
        .O(core__680_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__681
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[2]),
        .I4(core_n_272),
        .O(core__681_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__682
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(_T_2770[0]),
        .I4(core_n_271),
        .O(core__682_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__683
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(core_n_1687),
        .I4(core_n_270),
        .O(core__683_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__684
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(core_n_1686),
        .I4(core_n_269),
        .O(core__684_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__685
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(core_n_1685),
        .I4(core_n_268),
        .O(core__685_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__686
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(core_n_1684),
        .I4(core_n_267),
        .O(core__686_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__687
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(core_n_1683),
        .I4(core_n_266),
        .O(core__687_n_0));
  LUT5 #(
    .INIT(32'h0000FEEE)) 
    core__688
       (.I0(core_n_103),
        .I1(core_n_238),
        .I2(core_n_0),
        .I3(core_n_1682),
        .I4(core_n_265),
        .O(core__688_n_0));
  LUT6 #(
    .INIT(64'hF0D0F0F0F0D0D0D0)) 
    core__689
       (.I0(id_ctrl_rxs2),
        .I1(_T_1844),
        .I2(core__706_n_0),
        .I3(_GEN_274[1]),
        .I4(core_n_1249),
        .I5(_T_1416[1]),
        .O(ex_reg_rs_lsb_1[1]));
  LUT6 #(
    .INIT(64'h00000004FFFFFFFF)) 
    core__69
       (.I0(frontend_n_268),
        .I1(frontend_n_269),
        .I2(ibuf_io_inst_0_bits_raw[14]),
        .I3(ibuf_io_inst_0_bits_raw[0]),
        .I4(ibuf_io_inst_0_bits_raw[15]),
        .I5(ibuf_io_inst_0_bits_raw[1]),
        .O(core__69_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFDDFDD)) 
    core__690
       (.I0(id_ctrl_rxs2),
        .I1(_T_1844),
        .I2(core_n_1249),
        .I3(_T_1416[0]),
        .I4(_GEN_274[0]),
        .I5(core__705_n_0),
        .O(ex_reg_rs_lsb_1[0]));
  LUT3 #(
    .INIT(8'h20)) 
    core__691
       (.I0(id_ctrl_rxs2),
        .I1(_T_1844),
        .I2(_T_1790),
        .O(core__691_n_0));
  LUT6 #(
    .INIT(64'hFD20FFFFFD200000)) 
    core__692
       (.I0(frontend_n_388),
        .I1(_T_1829),
        .I2(core_n_1129),
        .I3(core__49_n_0),
        .I4(frontend_n_352),
        .I5(ibuf_io_inst_0_bits_raw[1]),
        .O(core__692_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2499" *) 
  LUT4 #(
    .INIT(16'h20F0)) 
    core__693
       (.I0(frontend_n_388),
        .I1(_T_1829),
        .I2(_T_1790),
        .I3(frontend_n_352),
        .O(ex_reg_rs_msb_0));
  LUT6 #(
    .INIT(64'h035703FFFFFFFFFF)) 
    core__694
       (.I0(_T_1031[14]),
        .I1(_T_1031[3]),
        .I2(_T_1005[4]),
        .I3(_T_1050[2]),
        .I4(_T_1005[6]),
        .I5(frontend_n_390),
        .O(id_ctrl_sel_alu1[0]));
  (* SOFT_HLUTNM = "soft_lutpair2495" *) 
  LUT4 #(
    .INIT(16'hFFF7)) 
    core__695
       (.I0(_T_1142[13]),
        .I1(_T_1031[3]),
        .I2(_T_1031[14]),
        .I3(_T_1005[6]),
        .O(core__695_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2544" *) 
  LUT3 #(
    .INIT(8'h80)) 
    core__696
       (.I0(_T_1142[13]),
        .I1(_T_1031[3]),
        .I2(frontend_n_366),
        .O(id_ctrl_mem_cmd[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    core__697
       (.I0(_T_889[24]),
        .I1(_T_877),
        .I2(frontend_n_402),
        .I3(frontend_n_226),
        .I4(_T_889[22]),
        .I5(_T_889[21]),
        .O(core__697_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2486" *) 
  LUT5 #(
    .INIT(32'h04440404)) 
    core__698
       (.I0(_T_1050[2]),
        .I1(_T_1005[4]),
        .I2(_T_1005[6]),
        .I3(_T_1050[5]),
        .I4(_T_1142[13]),
        .O(core__698_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2486" *) 
  LUT3 #(
    .INIT(8'h10)) 
    core__699
       (.I0(_T_1005[4]),
        .I1(_T_1050[2]),
        .I2(_T_1005[6]),
        .O(core__699_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__7
       (.I0(_GEN_274[63]),
        .I1(frontend_n_351),
        .I2(_T_1406[63]),
        .I3(frontend_n_352),
        .O(core__7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2482" *) 
  LUT5 #(
    .INIT(32'h00000100)) 
    core__70
       (.I0(ibuf_io_inst_0_bits_raw[15]),
        .I1(ibuf_io_inst_0_bits_raw[0]),
        .I2(ibuf_io_inst_0_bits_raw[14]),
        .I3(frontend_n_269),
        .I4(frontend_n_268),
        .O(core__70_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2481" *) 
  LUT4 #(
    .INIT(16'h44F4)) 
    core__700
       (.I0(_T_1005[4]),
        .I1(_T_1031[3]),
        .I2(_T_1005[6]),
        .I3(_T_1050[2]),
        .O(id_ctrl_sel_imm[0]));
  (* SOFT_HLUTNM = "soft_lutpair2493" *) 
  LUT4 #(
    .INIT(16'h44F4)) 
    core__701
       (.I0(_T_1005[4]),
        .I1(_T_1031[3]),
        .I2(_T_1050[2]),
        .I3(_T_1005[6]),
        .O(id_ctrl_sel_imm[1]));
  (* SOFT_HLUTNM = "soft_lutpair2481" *) 
  LUT5 #(
    .INIT(32'hFFFBFFFF)) 
    core__702
       (.I0(_T_1005[4]),
        .I1(_T_1031[3]),
        .I2(_T_1050[5]),
        .I3(_T_1005[6]),
        .I4(_T_1050[2]),
        .O(core__702_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2493" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    core__703
       (.I0(_T_1005[4]),
        .I1(_T_1031[3]),
        .I2(_T_1005[6]),
        .I3(frontend_n_396),
        .O(id_ctrl_fence_i));
  LUT6 #(
    .INIT(64'hFF0FFF0FFF0FBB0B)) 
    core__704
       (.I0(_T_1005[4]),
        .I1(_T_1031[3]),
        .I2(_T_909[26]),
        .I3(core__695_n_0),
        .I4(frontend_n_364),
        .I5(_T_1005[6]),
        .O(core__704_n_0));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FFF7)) 
    core__705
       (.I0(ex_ctrl_wxd),
        .I1(ex_reg_valid),
        .I2(frontend_n_375),
        .I3(frontend_n_362),
        .I4(mem_ctrl_mem),
        .I5(core_n_1093),
        .O(core__705_n_0));
  LUT4 #(
    .INIT(16'h00F7)) 
    core__706
       (.I0(ex_ctrl_wxd),
        .I1(ex_reg_valid),
        .I2(frontend_n_375),
        .I3(frontend_n_362),
        .O(core__706_n_0));
  LUT5 #(
    .INIT(32'h04040400)) 
    core__707
       (.I0(mem_reg_replay_reg),
        .I1(ex_reg_valid),
        .I2(core_n_1317),
        .I3(ex_reg_xcpt),
        .I4(ex_reg_xcpt_interrupt),
        .O(mem_reg_xcpt0));
  LUT5 #(
    .INIT(32'hFFF10001)) 
    core__708
       (.I0(core_n_1320),
        .I1(core__201_n_0),
        .I2(mem_reg_xcpt_interrupt),
        .I3(mem_reg_xcpt),
        .I4(mem_reg_cause[2]),
        .O(core__708_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    core__708_i_12
       (.I0(csr_io_bp_0_address[38]),
        .I1(core_n_1329),
        .O(core__708_i_12_n_0));
  CARRY4 core__708_i_16
       (.CI(core__708_i_30_n_0),
        .CO({core__708_i_16_n_0,core__708_i_16_n_1,core__708_i_16_n_2,core__708_i_16_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_2155,core_n_2156,core_n_2157,core_n_2158}));
  CARRY4 core__708_i_21
       (.CI(core__708_i_35_n_0),
        .CO({core__708_i_21_n_0,core__708_i_21_n_1,core__708_i_21_n_2,core__708_i_21_n_3}),
        .CYINIT(\<const0> ),
        .DI({core_n_2184,core_n_2185,core_n_2186,core_n_2187}),
        .S({core_n_2180,core_n_2181,core_n_2182,core_n_2183}));
  CARRY4 core__708_i_30
       (.CI(\<const0> ),
        .CO({core__708_i_30_n_0,core__708_i_30_n_1,core__708_i_30_n_2,core__708_i_30_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_2151,core_n_2152,core_n_2153,core_n_2154}));
  CARRY4 core__708_i_35
       (.CI(core__708_i_48_n_0),
        .CO({core__708_i_35_n_0,core__708_i_35_n_1,core__708_i_35_n_2,core__708_i_35_n_3}),
        .CYINIT(\<const0> ),
        .DI({core_n_2176,core_n_2177,core_n_2178,core_n_2179}),
        .S({core_n_2172,core_n_2173,core_n_2174,core_n_2175}));
  CARRY4 core__708_i_4
       (.CI(core__708_i_6_n_0),
        .CO(\bpu/_T_66 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,core_n_2163}));
  CARRY4 core__708_i_48
       (.CI(\<const0> ),
        .CO({core__708_i_48_n_0,core__708_i_48_n_1,core__708_i_48_n_2,core__708_i_48_n_3}),
        .CYINIT(\<const1> ),
        .DI({core_n_2168,core_n_2169,core_n_2170,core_n_2171}),
        .S({core_n_2164,core_n_2165,core_n_2166,core_n_2167}));
  CARRY4 core__708_i_5
       (.CI(core__708_i_8_n_0),
        .CO({\bpu/_T_39 ,core__708_i_5_n_1,core__708_i_5_n_2,core__708_i_5_n_3}),
        .CYINIT(\<const0> ),
        .DI({core__323_n_0,core_n_2199,core_n_2200,core_n_2201}),
        .S({core__708_i_12_n_0,core_n_2196,core_n_2197,core_n_2198}));
  CARRY4 core__708_i_6
       (.CI(core__708_i_16_n_0),
        .CO({core__708_i_6_n_0,core__708_i_6_n_1,core__708_i_6_n_2,core__708_i_6_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_2159,core_n_2160,core_n_2161,core_n_2162}));
  CARRY4 core__708_i_8
       (.CI(core__708_i_21_n_0),
        .CO({core__708_i_8_n_0,core__708_i_8_n_1,core__708_i_8_n_2,core__708_i_8_n_3}),
        .CYINIT(\<const0> ),
        .DI({core_n_2192,core_n_2193,core_n_2194,core_n_2195}),
        .S({core_n_2188,core_n_2189,core_n_2190,core_n_2191}));
  LUT5 #(
    .INIT(32'hFFF10001)) 
    core__709
       (.I0(core_n_1320),
        .I1(core__201_n_0),
        .I2(mem_reg_xcpt_interrupt),
        .I3(mem_reg_xcpt),
        .I4(mem_reg_cause[3]),
        .O(core__709_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2477" *) 
  LUT5 #(
    .INIT(32'h11111011)) 
    core__71
       (.I0(ibuf_io_inst_0_bits_raw[0]),
        .I1(ibuf_io_inst_0_bits_raw[1]),
        .I2(ibuf_io_inst_0_bits_raw[14]),
        .I3(frontend_n_269),
        .I4(ibuf_io_inst_0_bits_raw[15]),
        .O(core__71_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2484" *) 
  LUT5 #(
    .INIT(32'hFDFFFD00)) 
    core__710
       (.I0(mem_ctrl_branch),
        .I1(core_n_1345),
        .I2(core_n_1346),
        .I3(core_n_1347),
        .I4(core_n_1348),
        .O(core__710_n_0));
  LUT5 #(
    .INIT(32'hC55FC550)) 
    core__711
       (.I0(core_n_1775),
        .I1(mem_reg_rs2[41]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[1]),
        .O(mem_reg_rs20_in[41]));
  LUT6 #(
    .INIT(64'hCFC05F5FCFC05050)) 
    core__712
       (.I0(core_n_1775),
        .I1(mem_reg_rs2[57]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[25]),
        .I4(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I5(mem_reg_rs2[1]),
        .O(mem_reg_rs20_in[57]));
  LUT3 #(
    .INIT(8'hC5)) 
    core__713
       (.I0(core_n_1775),
        .I1(\div/_T_94 ),
        .I2(core_n_103),
        .O(\div/p_1_in ));
  LUT4 #(
    .INIT(16'hFF04)) 
    core__714
       (.I0(frontend_n_364),
        .I1(frontend_n_367),
        .I2(frontend_n_226),
        .I3(frontend_n_361),
        .O(core__714_n_0));
  LUT6 #(
    .INIT(64'hFFFF0404FF00FF00)) 
    core__715
       (.I0(frontend_n_364),
        .I1(frontend_n_367),
        .I2(frontend_n_226),
        .I3(core_n_91),
        .I4(frontend_n_230),
        .I5(_T_1790),
        .O(core__715_n_0));
  LUT5 #(
    .INIT(32'h10101000)) 
    core__716
       (.I0(core_n_101),
        .I1(target_reset),
        .I2(core_n_103),
        .I3(core_n_104),
        .I4(core_n_98),
        .O(core__716_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    core__717
       (.I0(\fq/elts_0_pc ),
        .I1(frontend_n_54),
        .I2(s2_pc[38]),
        .I3(\ibuf/_T_100 ),
        .I4(core_n_1070),
        .I5(csr_io_bp_0_address[38]),
        .O(core__717_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2553" *) 
  LUT3 #(
    .INIT(8'hAE)) 
    core__72
       (.I0(ibuf_io_inst_0_bits_raw[15]),
        .I1(frontend_n_269),
        .I2(ibuf_io_inst_0_bits_raw[14]),
        .O(core__72_n_0));
  LUT6 #(
    .INIT(64'hFBF80B08FFFFFFFF)) 
    core__73
       (.I0(frontend_io_cpu_resp_bits_data[30]),
        .I1(frontend_io_cpu_resp_bits_pc[1]),
        .I2(\ibuf/_T_100 ),
        .I3(frontend_io_cpu_resp_bits_data[14]),
        .I4(core_n_2087),
        .I5(frontend_n_269),
        .O(core__73_n_0));
  LUT4 #(
    .INIT(16'h4555)) 
    core__74
       (.I0(ibuf_io_inst_0_bits_raw[5]),
        .I1(frontend_n_268),
        .I2(ibuf_io_inst_0_bits_raw[11]),
        .I3(frontend_n_269),
        .O(core__74_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2480" *) 
  LUT5 #(
    .INIT(32'h0001FFFF)) 
    core__75
       (.I0(ibuf_io_inst_0_bits_raw[15]),
        .I1(ibuf_io_inst_0_bits_raw[0]),
        .I2(ibuf_io_inst_0_bits_raw[1]),
        .I3(frontend_n_269),
        .I4(ibuf_io_inst_0_bits_raw[6]),
        .O(core__75_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2477" *) 
  LUT5 #(
    .INIT(32'h00C40000)) 
    core__76
       (.I0(frontend_n_269),
        .I1(ibuf_io_inst_0_bits_raw[15]),
        .I2(ibuf_io_inst_0_bits_raw[14]),
        .I3(ibuf_io_inst_0_bits_raw[0]),
        .I4(ibuf_io_inst_0_bits_raw[1]),
        .O(core__76_n_0));
  LUT6 #(
    .INIT(64'h0407F4F7FFFFFFFF)) 
    core__77
       (.I0(frontend_io_cpu_resp_bits_data[29]),
        .I1(frontend_io_cpu_resp_bits_pc[1]),
        .I2(\ibuf/_T_100 ),
        .I3(frontend_io_cpu_resp_bits_data[13]),
        .I4(core_n_2088),
        .I5(ibuf_io_inst_0_bits_raw[15]),
        .O(core__77_n_0));
  LUT6 #(
    .INIT(64'h0000000D0000FF0D)) 
    core__78
       (.I0(ibuf_io_inst_0_bits_raw[14]),
        .I1(frontend_n_269),
        .I2(frontend_n_267),
        .I3(ibuf_io_inst_0_bits_raw[15]),
        .I4(ibuf_io_inst_0_bits_raw[1]),
        .I5(ibuf_io_inst_0_bits_raw[0]),
        .O(core__78_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    core__79
       (.I0(ibuf_io_inst_0_bits_raw[14]),
        .I1(ibuf_io_inst_0_bits_raw[3]),
        .I2(ibuf_io_inst_0_bits_raw[4]),
        .I3(ibuf_io_inst_0_bits_raw[2]),
        .I4(ibuf_io_inst_0_bits_raw[5]),
        .I5(ibuf_io_inst_0_bits_raw[6]),
        .O(core__79_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__8
       (.I0(_GEN_274[62]),
        .I1(frontend_n_351),
        .I2(_T_1406[62]),
        .I3(frontend_n_352),
        .O(core__8_n_0));
  LUT5 #(
    .INIT(32'h00000001)) 
    core__80
       (.I0(ibuf_io_inst_0_bits_raw[6]),
        .I1(ibuf_io_inst_0_bits_raw[5]),
        .I2(ibuf_io_inst_0_bits_raw[2]),
        .I3(ibuf_io_inst_0_bits_raw[4]),
        .I4(ibuf_io_inst_0_bits_raw[3]),
        .O(core__80_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2488" *) 
  LUT5 #(
    .INIT(32'hEF00FFFF)) 
    core__81
       (.I0(ibuf_io_inst_0_bits_raw[3]),
        .I1(ibuf_io_inst_0_bits_raw[1]),
        .I2(ibuf_io_inst_0_bits_raw[14]),
        .I3(ibuf_io_inst_0_bits_raw[0]),
        .I4(ibuf_io_inst_0_bits_raw[15]),
        .O(core__81_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2494" *) 
  LUT4 #(
    .INIT(16'h1000)) 
    core__82
       (.I0(ibuf_io_inst_0_bits_raw[1]),
        .I1(frontend_n_267),
        .I2(ibuf_io_inst_0_bits_raw[15]),
        .I3(ibuf_io_inst_0_bits_raw[14]),
        .O(core__82_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2500" *) 
  LUT4 #(
    .INIT(16'h0100)) 
    core__83
       (.I0(ibuf_io_inst_0_bits_raw[1]),
        .I1(frontend_n_267),
        .I2(ibuf_io_inst_0_bits_raw[15]),
        .I3(ibuf_io_inst_0_bits_raw[14]),
        .O(core__83_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2494" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    core__84
       (.I0(ibuf_io_inst_0_bits_raw[14]),
        .I1(ibuf_io_inst_0_bits_raw[1]),
        .I2(frontend_n_267),
        .I3(ibuf_io_inst_0_bits_raw[15]),
        .O(core__84_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2488" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    core__85
       (.I0(ibuf_io_inst_0_bits_raw[0]),
        .I1(ibuf_io_inst_0_bits_raw[1]),
        .I2(ibuf_io_inst_0_bits_raw[15]),
        .O(core__85_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2480" *) 
  LUT3 #(
    .INIT(8'h40)) 
    core__86
       (.I0(ibuf_io_inst_0_bits_raw[0]),
        .I1(ibuf_io_inst_0_bits_raw[1]),
        .I2(ibuf_io_inst_0_bits_raw[15]),
        .O(core__86_n_0));
  LUT6 #(
    .INIT(64'hFFEFFFEAAAEFAAEA)) 
    core__87
       (.I0(ibuf_io_inst_0_bits_raw[15]),
        .I1(frontend_io_cpu_resp_bits_data[26]),
        .I2(frontend_io_cpu_resp_bits_pc[1]),
        .I3(\ibuf/_T_100 ),
        .I4(frontend_io_cpu_resp_bits_data[10]),
        .I5(core_n_2091),
        .O(core__87_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2500" *) 
  LUT3 #(
    .INIT(8'h01)) 
    core__88
       (.I0(ibuf_io_inst_0_bits_raw[15]),
        .I1(frontend_n_267),
        .I2(ibuf_io_inst_0_bits_raw[1]),
        .O(core__88_n_0));
  LUT3 #(
    .INIT(8'hE0)) 
    core__89
       (.I0(ibuf_io_inst_0_bits_raw[15]),
        .I1(ibuf_io_inst_0_bits_raw[0]),
        .I2(ibuf_io_inst_0_bits_raw[1]),
        .O(core__89_n_0));
  LUT4 #(
    .INIT(16'hE200)) 
    core__9
       (.I0(_GEN_274[61]),
        .I1(frontend_n_351),
        .I2(_T_1406[61]),
        .I3(frontend_n_352),
        .O(core__9_n_0));
  (* SOFT_HLUTNM = "soft_lutpair2553" *) 
  LUT3 #(
    .INIT(8'h45)) 
    core__90
       (.I0(ibuf_io_inst_0_bits_raw[1]),
        .I1(frontend_n_267),
        .I2(ibuf_io_inst_0_bits_raw[15]),
        .O(core__90_n_0));
  LUT6 #(
    .INIT(64'hFB080000FFFFFFFF)) 
    core__91
       (.I0(frontend_io_cpu_resp_bits_data[3]),
        .I1(\ibuf/_T_100 ),
        .I2(frontend_io_cpu_resp_bits_pc[1]),
        .I3(frontend_io_cpu_resp_bits_data[19]),
        .I4(ibuf_io_inst_0_bits_raw[0]),
        .I5(ibuf_io_inst_0_bits_raw[1]),
        .O(core__91_n_0));
  LUT6 #(
    .INIT(64'h4044404040004040)) 
    core__92
       (.I0(frontend_n_267),
        .I1(ibuf_io_inst_0_bits_raw[1]),
        .I2(frontend_io_cpu_resp_bits_data[19]),
        .I3(frontend_io_cpu_resp_bits_pc[1]),
        .I4(\ibuf/_T_100 ),
        .I5(frontend_io_cpu_resp_bits_data[3]),
        .O(core__92_n_0));
  LUT4 #(
    .INIT(16'h6900)) 
    core__93
       (.I0(\ibuf/_T_100 ),
        .I1(frontend_n_265),
        .I2(frontend_io_cpu_resp_bits_pc[1]),
        .I3(frontend_io_cpu_resp_valid),
        .O(core__93_n_0));
  LUT6 #(
    .INIT(64'h55555555F7F5F7FF)) 
    core__94
       (.I0(frontend_n_265),
        .I1(core_n_68),
        .I2(frontend_io_ptw_status_prv[1]),
        .I3(ibuf_io_inst_0_bits_raw[25]),
        .I4(frontend_n_223),
        .I5(core_n_891),
        .O(core__94_n_0));
  LUT6 #(
    .INIT(64'h4540554045404540)) 
    core__95
       (.I0(core__128_n_0),
        .I1(core_n_95),
        .I2(\ibuf/_T_100 ),
        .I3(frontend_io_cpu_resp_bits_xcpt_pf_inst),
        .I4(ibuf_io_inst_0_bits_xcpt0_ae_inst),
        .I5(frontend_n_265),
        .O(core__95_n_0));
  LUT6 #(
    .INIT(64'h0000101000051015)) 
    core__96
       (.I0(core__128_n_0),
        .I1(core_n_95),
        .I2(\ibuf/_T_100 ),
        .I3(frontend_io_cpu_resp_bits_xcpt_pf_inst),
        .I4(\ibuf/buf__xcpt_ae_inst ),
        .I5(frontend_io_cpu_resp_bits_xcpt_ae_inst),
        .O(core__96_n_0));
  LUT6 #(
    .INIT(64'h5545004000000000)) 
    core__97
       (.I0(frontend_n_224),
        .I1(frontend_io_cpu_resp_bits_data[7]),
        .I2(\ibuf/_T_100 ),
        .I3(frontend_io_cpu_resp_bits_pc[1]),
        .I4(frontend_io_cpu_resp_bits_data[23]),
        .I5(ibuf_io_inst_0_bits_raw[22]),
        .O(core__97_n_0));
  LUT6 #(
    .INIT(64'h0000000000105515)) 
    core__98
       (.I0(ibuf_io_inst_0_bits_raw[22]),
        .I1(frontend_io_cpu_resp_bits_data[7]),
        .I2(\ibuf/_T_100 ),
        .I3(frontend_io_cpu_resp_bits_pc[1]),
        .I4(frontend_io_cpu_resp_bits_data[23]),
        .I5(frontend_n_224),
        .O(core__98_n_0));
  LUT6 #(
    .INIT(64'h0000457545754575)) 
    core__99
       (.I0(frontend_io_cpu_resp_bits_data[23]),
        .I1(frontend_io_cpu_resp_bits_pc[1]),
        .I2(\ibuf/_T_100 ),
        .I3(frontend_io_cpu_resp_bits_data[7]),
        .I4(frontend_n_224),
        .I5(frontend_n_222),
        .O(core__99_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep
       (.I0(alu_io_in1[1]),
        .I1(alu_io_in2[1]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__0
       (.I0(alu_io_in1[2]),
        .I1(alu_io_in2[2]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__0_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__1
       (.I0(alu_io_in1[3]),
        .I1(alu_io_in2[3]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__1_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__10
       (.I0(alu_io_in1[24]),
        .I1(alu_io_in2[24]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__10_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__11
       (.I0(alu_io_in1[27]),
        .I1(alu_io_in2[27]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__11_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__12
       (.I0(alu_io_in1[30]),
        .I1(alu_io_in2[30]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__12_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__13
       (.I0(alu_io_in1[33]),
        .I1(alu_io_in2[33]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__13_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__14
       (.I0(alu_io_in1[36]),
        .I1(alu_io_in2[36]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__14_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__15
       (.I0(alu_io_in1[39]),
        .I1(alu_io_in2[39]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__15_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__16
       (.I0(alu_io_in1[42]),
        .I1(alu_io_in2[42]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__16_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__17
       (.I0(alu_io_in1[45]),
        .I1(alu_io_in2[45]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__17_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__18
       (.I0(alu_io_in1[48]),
        .I1(alu_io_in2[48]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__18_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__19
       (.I0(alu_io_in1[51]),
        .I1(alu_io_in2[51]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__19_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__2
       (.I0(alu_io_in1[4]),
        .I1(alu_io_in2[4]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__2_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__20
       (.I0(alu_io_in1[54]),
        .I1(alu_io_in2[54]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__20_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__21
       (.I0(alu_io_in1[57]),
        .I1(alu_io_in2[57]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__21_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__22
       (.I0(alu_io_in1[60]),
        .I1(alu_io_in2[60]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__22_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core_rep__23
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core_rep__23_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core_rep__24
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core_rep__24_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core_rep__25
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core_rep__25_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core_rep__26
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core_rep__26_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core_rep__27
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core_rep__27_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core_rep__28
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core_rep__28_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core_rep__29
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core_rep__29_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__3
       (.I0(alu_io_in1[5]),
        .I1(alu_io_in2[5]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__3_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core_rep__30
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core_rep__30_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core_rep__31
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core_rep__31_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core_rep__32
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core_rep__32_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    core_rep__33
       (.I0(core_n_357),
        .I1(core_n_374),
        .O(core_rep__33_n_0));
  LUT4 #(
    .INIT(16'hAA8A)) 
    core_rep__34
       (.I0(core_n_1557),
        .I1(core_n_1347),
        .I2(core_n_1345),
        .I3(core_n_1346),
        .O(core_rep__34_n_0));
  LUT4 #(
    .INIT(16'h4404)) 
    core_rep__35
       (.I0(core_n_1013),
        .I1(core_n_1010),
        .I2(wb_reg_xcpt),
        .I3(wb_reg_cause),
        .O(core_rep__35_n_0));
  LUT4 #(
    .INIT(16'h0051)) 
    core_rep__36
       (.I0(core_n_1013),
        .I1(wb_reg_xcpt),
        .I2(wb_reg_cause),
        .I3(core_n_1010),
        .O(core_rep__36_n_0));
  LUT6 #(
    .INIT(64'h65AA65659A559A9A)) 
    core_rep__4
       (.I0(alu_io_in1[6]),
        .I1(core_n_1777),
        .I2(mem_reg_rs2[6]),
        .I3(core_n_1776),
        .I4(core_n_1243),
        .I5(ex_ctrl_alu_fn),
        .O(core_rep__4_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__5
       (.I0(alu_io_in1[11]),
        .I1(alu_io_in2[11]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__5_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__6
       (.I0(alu_io_in1[12]),
        .I1(alu_io_in2[12]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__6_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__7
       (.I0(alu_io_in1[15]),
        .I1(alu_io_in2[15]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__7_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__8
       (.I0(alu_io_in1[18]),
        .I1(alu_io_in2[18]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__8_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    core_rep__9
       (.I0(alu_io_in1[21]),
        .I1(alu_io_in2[21]),
        .I2(ex_ctrl_alu_fn),
        .O(core_rep__9_n_0));
  DCache dcache
       (.ADDRARDADDR(ADDRARDADDR),
        .CO(_T_2437),
        .D({_T_273,dcache_io_cpu_req_bits_addr[5:3],ptw_n_49,ptw_n_50,ptw_n_51}),
        .DIA(tlMasterXbar_auto_out_c_bits_size),
        .DIB({dcache_n_137,dcache_n_138}),
        .DOA(tlMasterXbar_auto_in_0_d_bits_opcode),
        .DOBDO({dcache_n_0,dcache_n_1,dcache_n_2,dcache_n_3,dcache_n_4,dcache_n_5,dcache_n_6,dcache_n_7}),
        .E(_T_258),
        .Q({dcache_n_139,dcache_n_140,dcache_n_141,dcache_n_142,dcache_n_143,dcache_n_144,dcache_n_145,dcache_n_146,dcache_n_147,dcache_n_148,dcache_n_149,dcache_n_150,dcache_n_151,dcache_n_152,dcache_n_153,dcache_n_154,dcache_n_155,dcache_n_156,dcache_n_157,dcache_n_158,dcache_n_159,_T_628}),
        .S({core_n_1994,ptw_n_190,core_n_1995,core_n_1996}),
        .\_T_1052_reg[2] (dcache_n_343),
        .\_T_1052_reg[3] (dcache_n_342),
        .\_T_1052_reg[7] (dcache_n_213),
        .\_T_1066_reg[1] (dcache_n_209),
        .\_T_1066_reg[1]_0 (tlMasterXbar_n_6),
        ._T_1161_0_reg(tlMasterXbar_n_10),
        ._T_1172_1(_T_1172_1),
        ._T_1208({_T_1208[114:110],_T_1208[106],_T_1208[104],_T_1208[77:72],_T_1208[63:0]}),
        ._T_1498(_T_1498),
        .\_T_1643_reg[7]_0 (tlMasterXbar_auto_out_c_bits_data),
        ._T_165_reg(frontend_n_49),
        ._T_1701(_T_1701),
        ._T_177(_T_177),
        ._T_179(_T_179),
        .\_T_1883_reg[0] (core_n_2079),
        .\_T_1883_reg[1] (core_n_1837),
        .\_T_1883_reg[1]_0 (core_n_1839),
        .\_T_1883_reg[1]_1 (dcache_io_ptw_status_dprv),
        .\_T_1883_reg[1]_2 (core_n_1841),
        .\_T_250_0_bits_mask_reg[7] (dcache_n_455),
        .\_T_250_0_bits_mask_reg[7]_0 (dcache_n_456),
        .\_T_2547_reg[1] (dcache_n_552),
        .\_T_2547_reg[1]_0 (dcache_n_553),
        .\_T_2547_reg[24] (dcache_n_550),
        .\_T_2547_reg[24]_0 (dcache_n_559),
        .\_T_2547_reg[25] (dcache_n_561),
        .\_T_2547_reg[26] (dcache_n_563),
        .\_T_2547_reg[27] (dcache_n_565),
        .\_T_2547_reg[28] (dcache_n_560),
        .\_T_2547_reg[29] (dcache_n_562),
        .\_T_2547_reg[30] (dcache_n_564),
        .\_T_2547_reg[30]_0 (core_n_1096),
        .\_T_2547_reg[31] (dcache_n_566),
        ._T_255(_T_255),
        .\_T_277_reg[2] (dcache_n_555),
        .\_T_281_reg[0] (dcache_n_556),
        .\_T_3585_reg[0]_0 (sync_xing_n_210),
        .\_T_3585_reg[0]_1 (p_0_in_5),
        .\_T_3585_reg[1]_0 (_T_3585_reg__0),
        .\_T_3585_reg[6]_0 (dcache_n_453),
        .\_T_3585_reg[8]_0 (dcache_n_212),
        .\_T_3585_reg[8]_1 (dcache_n_431),
        .\_T_3585_reg[8]_2 (dcache_n_432),
        ._T_3628(_T_3628),
        ._T_384(_T_384),
        .\_T_3859_reg[8]_0 (dcache_n_433),
        .\_T_386_reg[0] (ptw_n_82),
        .\_T_386_reg[0]_0 (ptw_n_83),
        .\_T_386_reg[2] (ptw_n_76),
        .\_T_389_reg[7] (_T_439),
        ._T_4068_pf_ld_reg_0(dcache_n_134),
        ._T_4068_pf_ld_reg_1({\tlb/entries_2_u ,\tlb/entries_2_sx ,\tlb/entries_2_sr }),
        ._T_4068_pf_ld_reg_2({\tlb/entries_3_u ,\tlb/entries_3_sx ,\tlb/entries_3_sr }),
        ._T_4068_pf_ld_reg_3(\tlb/_GEN_36 ),
        ._T_4068_pf_st_reg_0(dcache_n_133),
        ._T_4068_pf_st_reg_1(\tlb/entries_1_u ),
        .\_T_407_0_reg[19] (dcache_n_571),
        ._T_407_1(_T_407_1),
        .\_T_407_1_reg[0] (dcache_n_368),
        .\_T_407_1_reg[10] (dcache_n_379),
        .\_T_407_1_reg[11] (dcache_n_380),
        .\_T_407_1_reg[12] (dcache_n_381),
        .\_T_407_1_reg[13] (dcache_n_382),
        .\_T_407_1_reg[14] (dcache_n_383),
        .\_T_407_1_reg[15] (dcache_n_384),
        .\_T_407_1_reg[16] (dcache_n_385),
        .\_T_407_1_reg[17] (dcache_n_386),
        .\_T_407_1_reg[18] (dcache_n_387),
        .\_T_407_1_reg[19] (dcache_n_388),
        .\_T_407_1_reg[19]_0 (dcache_n_567),
        .\_T_407_1_reg[1] (dcache_n_370),
        .\_T_407_1_reg[2] (dcache_n_371),
        .\_T_407_1_reg[3] (dcache_n_372),
        .\_T_407_1_reg[4] (dcache_n_373),
        .\_T_407_1_reg[5] (dcache_n_374),
        .\_T_407_1_reg[6] (dcache_n_375),
        .\_T_407_1_reg[7] (dcache_n_376),
        .\_T_407_1_reg[8] (dcache_n_377),
        .\_T_407_1_reg[9] (dcache_n_378),
        .\_T_407_2_reg[19] (dcache_n_569),
        .\_T_407_3_reg[19] (dcache_n_570),
        ._T_407_4(_T_407_4),
        .\_T_407_4_reg[19] (dcache_n_572),
        .\_T_407_5_reg[19] (dcache_n_573),
        ._T_407_6(_T_407_6),
        .\_T_407_6_reg[19] (dcache_n_574),
        .\_T_407_7_reg[19] (dcache_n_161),
        .\_T_407_7_reg[19]_0 (dcache_n_367),
        .\_T_407_7_reg[19]_1 (dcache_n_575),
        ._T_435(_T_435),
        ._T_481(_T_481),
        ._T_499(_T_499),
        .\_T_973_reg[1] (dcache_n_633),
        .blockProbeAfterGrantCount(blockProbeAfterGrantCount),
        .blockUncachedGrant(blockUncachedGrant),
        .blockUncachedGrant_reg_0(sync_xing_n_212),
        .blockUncachedGrant_reg_1(sync_xing_n_213),
        .blockUncachedGrant_reg_2(sync_xing_n_214),
        .blockUncachedGrant_reg_3(sync_xing_n_215),
        .blockUncachedGrant_reg_4(sync_xing_n_216),
        .blockUncachedGrant_reg_5(sync_xing_n_217),
        .blockUncachedGrant_reg_6(sync_xing_n_218),
        .buf__replay_reg(dcache_n_543),
        .buf__replay_reg_0(dcache_n_544),
        .\bypass_mux_2_reg[10] (core_n_1259),
        .\bypass_mux_2_reg[11] (core_n_1260),
        .\bypass_mux_2_reg[12] (core_n_1258),
        .\bypass_mux_2_reg[13] (core_n_1261),
        .\bypass_mux_2_reg[14] (core_n_1262),
        .\bypass_mux_2_reg[15] (core_n_1263),
        .\bypass_mux_2_reg[16] (core_n_1264),
        .\bypass_mux_2_reg[17] (core_n_1265),
        .\bypass_mux_2_reg[18] (core_n_1266),
        .\bypass_mux_2_reg[19] (core_n_1267),
        .\bypass_mux_2_reg[20] (core_n_1268),
        .\bypass_mux_2_reg[21] (core_n_1269),
        .\bypass_mux_2_reg[22] (core_n_1270),
        .\bypass_mux_2_reg[23] (core_n_1271),
        .\bypass_mux_2_reg[24] (core_n_1272),
        .\bypass_mux_2_reg[25] (core_n_1273),
        .\bypass_mux_2_reg[26] (core_n_1274),
        .\bypass_mux_2_reg[27] (core_n_1275),
        .\bypass_mux_2_reg[28] (core_n_1276),
        .\bypass_mux_2_reg[29] (core_n_1277),
        .\count_reg[1] (dcache_n_580),
        .\count_reg[1]_0 (ptw_n_37),
        .dataArb_io_in_1_bits_addr({dataArb_io_in_1_bits_addr[11],dataArb_io_in_1_bits_addr[9],dataArb_io_in_1_bits_addr[7:6]}),
        .dataArb_io_in_1_valid(dataArb_io_in_1_valid),
        .dataArb_io_in_2_valid(dataArb_io_in_2_valid),
        .data_arrays_0_0_reg(dcache_n_417),
        .data_arrays_0_0_reg_0(dcache_n_418),
        .data_arrays_0_0_reg_1(dcache_n_448),
        .data_arrays_0_0_reg_2(dcache_n_454),
        .data_arrays_0_0_reg_i_44(data_arrays_0_0_reg_i_44),
        .data_arrays_0_0_reg_i_45(data_arrays_0_0_reg_i_45),
        .data_arrays_0_0_reg_i_46(data_arrays_0_0_reg_i_46),
        .data_arrays_0_0_reg_i_47(data_arrays_0_0_reg_i_47),
        .data_arrays_0_0_reg_i_48(data_arrays_0_0_reg_i_48),
        .data_arrays_0_0_reg_i_49(data_arrays_0_0_reg_i_49),
        .data_arrays_0_0_reg_i_50(data_arrays_0_0_reg_i_50),
        .data_arrays_0_0_reg_i_51(data_arrays_0_0_reg_i_51),
        .data_arrays_0_0_reg_i_52(data_arrays_0_0_reg_i_52),
        .data_arrays_0_0_reg_i_52_0(data_arrays_0_0_reg_i_52_0),
        .data_arrays_0_7_reg(dcache_n_136),
        .data_arrays_0_7_reg_0(_T_766),
        .dcacheArb_io_requestor_0_req_ready(dcacheArb_io_requestor_0_req_ready),
        .dcacheArb_io_requestor_0_s1_kill(dcacheArb_io_requestor_0_s1_kill),
        .dcacheArb_io_requestor_1_ordered(dcacheArb_io_requestor_1_ordered),
        .dcacheArb_io_requestor_1_replay_next(dcacheArb_io_requestor_1_replay_next),
        .dcacheArb_io_requestor_1_req_bits_typ(dcacheArb_io_requestor_1_req_bits_typ),
        .dcacheArb_io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),
        .dcacheArb_io_requestor_1_resp_bits_data({dcacheArb_io_requestor_1_resp_bits_data[63:30],dcacheArb_io_requestor_1_resp_bits_data[9:0]}),
        .dcacheArb_io_requestor_1_resp_bits_data_word_bypass(dcacheArb_io_requestor_1_resp_bits_data_word_bypass),
        .dcacheArb_io_requestor_1_resp_bits_replay(dcacheArb_io_requestor_1_resp_bits_replay),
        .dcacheArb_io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),
        .dcacheArb_io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),
        .dcacheArb_io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),
        .dcacheArb_io_requestor_1_s2_xcpt_ae_ld(dcacheArb_io_requestor_1_s2_xcpt_ae_ld),
        .dcacheArb_io_requestor_1_s2_xcpt_ma_ld(dcacheArb_io_requestor_1_s2_xcpt_ma_ld),
        .dcacheArb_io_requestor_1_s2_xcpt_ma_st(dcacheArb_io_requestor_1_s2_xcpt_ma_st),
        .dcacheArb_io_requestor_1_s2_xcpt_pf_ld(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
        .dcacheArb_io_requestor_1_s2_xcpt_pf_st(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
        .dcache_io_cpu_invalidate_lr(dcache_io_cpu_invalidate_lr),
        .dcache_io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr[31:6]),
        .dcache_io_ptw_resp_bits_level(dcache_io_ptw_resp_bits_level),
        .dcache_io_ptw_resp_bits_pte_v(dcache_io_ptw_resp_bits_pte_v),
        .dcache_io_ptw_resp_valid(dcache_io_ptw_resp_valid),
        .dcache_io_ptw_status_mxr(dcache_io_ptw_status_mxr),
        .dcache_io_ptw_status_sum(dcache_io_ptw_status_sum),
        .doUncachedResp_reg_0(core_n_1095),
        .\ex_ctrl_mem_cmd_reg[4] (dcacheArb_io_requestor_1_req_bits_cmd),
        .\ex_ctrl_mem_cmd_reg[4]_0 (core_n_1028),
        .ex_ctrl_mem_reg(dcache_n_541),
        .ex_ctrl_mem_reg_0(dcache_n_542),
        .ex_ctrl_mem_reg_1(dcache_n_551),
        .\ex_reg_inst_reg[11] (dcacheArb_io_requestor_1_req_bits_tag),
        .\ex_reg_rs_msb_0_reg[27] (_GEN_274[29:10]),
        .\ex_reg_rs_msb_0_reg[8] (dcache_n_369),
        .\ex_reg_rs_msb_1_reg[61] (dcache_n_554),
        .frontend_io_ptw_pmp_1_cfg_a(frontend_io_ptw_pmp_1_cfg_a),
        .frontend_io_ptw_pmp_1_cfg_w(frontend_io_ptw_pmp_1_cfg_w),
        .frontend_io_ptw_pmp_2_cfg_a(frontend_io_ptw_pmp_2_cfg_a),
        .frontend_io_ptw_pmp_6_cfg_a(frontend_io_ptw_pmp_6_cfg_a),
        .frontend_io_ptw_pmp_7_cfg_a(frontend_io_ptw_pmp_7_cfg_a),
        .frontend_io_ptw_ptbr_mode(frontend_io_ptw_ptbr_mode),
        .grantInProgress_reg_0(dcache_n_75),
        .grantInProgress_reg_1(sync_xing_n_51),
        .host_clk(host_clk),
        .ibuf_io_inst_0_bits_inst_rd({ibuf_io_inst_0_bits_inst_rd[4],ibuf_io_inst_0_bits_inst_rd[1:0]}),
        .ibuf_io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
        .ibuf_io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
        .invalid_paddr(invalid_paddr),
        .io_enq_bits_address(tlMasterXbar_auto_out_c_bits_address),
        .io_enq_bits_mask(tlMasterXbar_auto_out_a_bits_mask[5:0]),
        .io_enq_bits_source(tlMasterXbar_auto_out_c_bits_source),
        .\lrscAddr_reg[25]_0 ({_GEN_283_0,_T_3959}),
        .\lrscCount_reg[4]_0 (dcache_n_435),
        .maybe_full(\Queue_3/maybe_full ),
        .maybe_full_reg(sync_xing_n_32),
        .maybe_full_reg_0(sync_xing_n_22),
        .\mem_reg_rs2_reg[63] (dcacheArb_io_requestor_1_s1_data_data),
        .nBufValid_reg(frontend_n_387),
        .pte_v(pte_v),
        .r_pte_a_reg(dcache_n_443),
        .r_pte_a_reg_0(dcache_n_583),
        .r_pte_d(r_pte_d),
        .r_pte_d_reg({\tlb/_T_936 ,\tlb/_T_943 ,\tlb/_T_928 ,\tlb/_T_949 ,\tlb/_T_946 }),
        .r_pte_g_reg(dcache_n_442),
        .\r_pte_ppn_reg[19] ({ptw_n_154,core_n_1875,core_n_1876}),
        .\r_pte_ppn_reg[19]_0 ({ptw_n_157,core_n_1877,core_n_1878}),
        .\r_pte_ppn_reg[19]_1 ({ptw_n_147,core_n_1873,core_n_1874}),
        .\r_pte_ppn_reg[19]_2 ({ptw_n_141,core_n_1869,core_n_1870}),
        .\r_pte_ppn_reg[19]_3 ({ptw_n_144,core_n_1871,core_n_1872}),
        .\r_pte_ppn_reg[19]_4 ({ptw_n_150,ptw_n_151,core_n_1868}),
        .\r_pte_ppn_reg[19]_5 (\tlb/_T_382_3 ),
        .\r_pte_ppn_reg[19]_6 (\tlb/_T_392 ),
        .\r_pte_ppn_reg[19]_7 (dcache_io_ptw_resp_bits_pte_ppn),
        .r_pte_r_reg(dcache_n_438),
        .r_pte_u_reg(dcache_n_441),
        .r_pte_u_reg_0({dcache_io_ptw_resp_bits_pte_u,dcache_io_ptw_resp_bits_pte_g,dcache_io_ptw_resp_bits_ae}),
        .r_pte_v_reg(dcache_n_582),
        .r_pte_w_reg(dcache_n_439),
        .r_pte_x_reg(dcache_n_440),
        .ram_address__T_63_data(tlMasterXbar_auto_in_0_b_bits_address),
        .ram_data__T_63_data(tlMasterXbar_auto_in_0_d_bits_data),
        .\ram_id_reg[0] (tlMasterXbar_auto_out_c_bits_opcode),
        .ram_param__T_63_data(tlMasterXbar_auto_in_0_b_bits_param),
        .\reg_entries_0_reg[0] (dcache_n_584),
        .\reg_entries_0_reg[0]_0 ({\tlb/p_0_in ,\tlb/entries_4_u ,\tlb/entries_4_sx ,\tlb/entries_4_sr }),
        .\reg_entries_0_reg[0]_1 ({dcache_n_610,dcache_n_611}),
        .\reg_entries_0_reg[0]_2 (dcache_n_612),
        .\reg_entries_0_reg[0]_3 (dcache_n_635),
        .\reg_entries_0_reg[0]_4 ({dcache_n_636,dcache_n_637}),
        .\reg_entries_0_reg[0]_5 (dcache_n_638),
        .\reg_entries_0_reg[0]_6 (dcache_n_639),
        .\reg_entries_0_reg[0]_7 (dcache_n_640),
        .\reg_entries_0_reg[0]_8 (dcache_n_641),
        .\reg_entries_0_reg[10] (core_n_1838),
        .\reg_entries_0_reg[1] (dcache_n_642),
        .\reg_entries_0_reg[2] (dcache_n_643),
        .\reg_entries_0_reg[41] (dcache_io_ptw_req_bits_addr),
        .\reg_entries_0_reg[4] (\tlb/pmp/_T_74 ),
        .\reg_entries_0_reg[4]_0 (\tlb/pmp/_T_94 ),
        .\reg_entries_0_reg[4]_1 (dcache_n_614),
        .\reg_entries_0_reg[4]_2 (dcache_n_615),
        .\reg_entries_0_reg[4]_3 (dcache_n_621),
        .\reg_entries_0_reg[4]_4 (dcache_n_627),
        .\reg_entries_0_reg[4]_5 (dcache_n_629),
        .\reg_entries_0_reg[4]_6 (dcache_n_630),
        .\reg_entries_0_reg[4]_7 (dcache_n_631),
        .\reg_entries_0_reg[4]_8 (dcache_n_632),
        .\reg_entries_0_reg[6] (\tlb/pmp/_T_201 ),
        .\reg_entries_0_reg[6]_0 (\tlb/pmp/_T_328 ),
        .\reg_entries_0_reg[6]_1 (\tlb/pmp/_T_455 ),
        .\reg_entries_0_reg[6]_10 (dcache_n_619),
        .\reg_entries_0_reg[6]_11 (dcache_n_620),
        .\reg_entries_0_reg[6]_12 (dcache_n_622),
        .\reg_entries_0_reg[6]_13 (dcache_n_623),
        .\reg_entries_0_reg[6]_14 (dcache_n_624),
        .\reg_entries_0_reg[6]_15 (dcache_n_625),
        .\reg_entries_0_reg[6]_16 (dcache_n_626),
        .\reg_entries_0_reg[6]_17 (dcache_n_628),
        .\reg_entries_0_reg[6]_2 (\tlb/pmp/_T_582 ),
        .\reg_entries_0_reg[6]_3 (\tlb/pmp/_T_709 ),
        .\reg_entries_0_reg[6]_4 (\tlb/pmp/_T_836 ),
        .\reg_entries_0_reg[6]_5 (dcache_n_585),
        .\reg_entries_0_reg[6]_6 (dcache_n_613),
        .\reg_entries_0_reg[6]_7 (dcache_n_616),
        .\reg_entries_0_reg[6]_8 (dcache_n_617),
        .\reg_entries_0_reg[6]_9 (dcache_n_618),
        .\reg_entries_4_reg[57] ({ptw_n_186,ptw_n_187}),
        .\reg_entries_4_reg[57]_0 (ptw_n_166),
        .\reg_entries_4_reg[57]_1 ({ptw_n_188,ptw_n_189}),
        .\reg_entries_4_reg[57]_2 (ptw_n_185),
        .\reg_entries_4_reg[61] (\tlb/_T_728 ),
        .\reg_entries_4_reg[61]_0 (\tlb/_T_482 ),
        .reg_mstatus_mxr_reg(core_n_2084),
        .reg_mstatus_mxr_reg_0(core_n_2082),
        .reg_mstatus_sum_reg(core_n_2083),
        .reg_mstatus_sum_reg_0(core_n_2081),
        .reg_mstatus_sum_reg_1(core_n_2080),
        .reg_mstatus_sum_reg_2(core_n_2085),
        .\reg_pmp_0_addr_reg[16] ({core_n_1947,core_n_1948,core_n_1949,core_n_1950}),
        .\reg_pmp_0_addr_reg[16]_0 ({core_n_1943,core_n_1944,core_n_1945,core_n_1946}),
        .\reg_pmp_0_addr_reg[24] ({core_n_1883,core_n_1884,core_n_1885,core_n_1886}),
        .\reg_pmp_0_addr_reg[24]_0 ({core_n_1879,core_n_1880,core_n_1881,core_n_1882}),
        .\reg_pmp_0_addr_reg[29] ({core_n_1865,core_n_1866,core_n_1867}),
        .\reg_pmp_0_addr_reg[29]_0 ({frontend_io_ptw_pmp_0_addr[29],frontend_io_ptw_pmp_0_addr[8:1]}),
        .\reg_pmp_0_addr_reg[8] ({core_n_2056,core_n_2057,core_n_2058,core_n_2059}),
        .\reg_pmp_0_addr_reg[8]_0 ({core_n_2052,core_n_2053,core_n_2054,core_n_2055}),
        .\reg_pmp_0_addr_reg[8]_1 (core_n_2060),
        .\reg_pmp_1_addr_reg[16] ({core_n_1951,core_n_1952,core_n_1953,core_n_1954}),
        .\reg_pmp_1_addr_reg[16]_0 ({core_n_1983,core_n_1984,core_n_1985,core_n_1986}),
        .\reg_pmp_1_addr_reg[23] ({core_n_1932,core_n_1933,core_n_1934,ptw_n_192}),
        .\reg_pmp_1_addr_reg[24] ({core_n_1903,core_n_1904,core_n_1905,core_n_1906}),
        .\reg_pmp_1_addr_reg[29] ({core_n_1862,core_n_1863,core_n_1864}),
        .\reg_pmp_1_addr_reg[29]_0 ({core_n_391,core_n_392,core_n_393}),
        .\reg_pmp_1_addr_reg[6] (core_n_2051),
        .\reg_pmp_1_addr_reg[7] ({core_n_2043,core_n_2044,core_n_2045,core_n_2046}),
        .\reg_pmp_1_addr_reg[8] ({core_n_2047,core_n_2048,core_n_2049,core_n_2050}),
        .\reg_pmp_1_addr_reg[8]_0 ({frontend_io_ptw_pmp_1_addr[8:7],frontend_io_ptw_pmp_1_addr[5:0]}),
        .reg_pmp_1_cfg_r_reg(core_n_1835),
        .\reg_pmp_2_addr_reg[0] (ptw_n_139),
        .\reg_pmp_2_addr_reg[11] (ptw_n_140),
        .\reg_pmp_2_addr_reg[16] ({core_n_1955,core_n_1956,core_n_1957,core_n_1958}),
        .\reg_pmp_2_addr_reg[16]_0 ({core_n_1987,core_n_1988,ptw_n_179,core_n_1989}),
        .\reg_pmp_2_addr_reg[23] ({core_n_1887,core_n_1888,core_n_1889,core_n_1890}),
        .\reg_pmp_2_addr_reg[24] ({core_n_1891,core_n_1892,core_n_1893,core_n_1894}),
        .\reg_pmp_2_addr_reg[29] ({core_n_1859,core_n_1860,core_n_1861}),
        .\reg_pmp_2_addr_reg[29]_0 ({core_n_424,core_n_425,core_n_426}),
        .\reg_pmp_2_addr_reg[29]_1 ({frontend_io_ptw_pmp_2_addr[29],frontend_io_ptw_pmp_2_addr[8:0]}),
        .\reg_pmp_2_addr_reg[6] (core_n_2042),
        .\reg_pmp_2_addr_reg[7] ({core_n_2038,core_n_2039,core_n_2040,core_n_2041}),
        .\reg_pmp_2_addr_reg[8] ({core_n_2034,core_n_2035,core_n_2036,core_n_2037}),
        .\reg_pmp_3_addr_reg[16] ({core_n_1959,core_n_1960,core_n_1961,core_n_1962}),
        .\reg_pmp_3_addr_reg[16]_0 ({core_n_1990,core_n_1991,core_n_1992,core_n_1993}),
        .\reg_pmp_3_addr_reg[23] ({core_n_1895,core_n_1896,core_n_1897,core_n_1898}),
        .\reg_pmp_3_addr_reg[24] ({core_n_1899,core_n_1900,core_n_1901,core_n_1902}),
        .\reg_pmp_3_addr_reg[29] ({core_n_1856,core_n_1857,core_n_1858}),
        .\reg_pmp_3_addr_reg[6] (core_n_2024),
        .\reg_pmp_3_addr_reg[7] ({core_n_2016,core_n_2017,core_n_2018,core_n_2019}),
        .\reg_pmp_3_addr_reg[8] ({core_n_2020,core_n_2021,core_n_2022,core_n_2023}),
        .\reg_pmp_3_addr_reg[8]_0 ({frontend_io_ptw_pmp_3_addr[8:7],frontend_io_ptw_pmp_3_addr[5:0]}),
        .\reg_pmp_4_addr_reg[0] (ptw_n_142),
        .\reg_pmp_4_addr_reg[16] ({core_n_1963,core_n_1964,core_n_1965,core_n_1966}),
        .\reg_pmp_4_addr_reg[16]_0 ({core_n_2000,ptw_n_175,core_n_2001,core_n_2002}),
        .\reg_pmp_4_addr_reg[24] ({core_n_1907,core_n_1908,core_n_1909,core_n_1910}),
        .\reg_pmp_4_addr_reg[24]_0 ({core_n_1939,core_n_1940,core_n_1941,core_n_1942}),
        .\reg_pmp_4_addr_reg[29] ({core_n_1853,core_n_1854,core_n_1855}),
        .\reg_pmp_4_addr_reg[29]_0 ({frontend_io_ptw_pmp_4_addr[29],frontend_io_ptw_pmp_4_addr[8:0]}),
        .\reg_pmp_4_addr_reg[4] (core_n_2015),
        .\reg_pmp_4_addr_reg[7] ({core_n_2011,core_n_2012,core_n_2013,core_n_2014}),
        .\reg_pmp_4_addr_reg[8] ({core_n_2007,core_n_2008,core_n_2009,core_n_2010}),
        .\reg_pmp_5_addr_reg[16] ({core_n_1967,core_n_1968,core_n_1969,core_n_1970}),
        .\reg_pmp_5_addr_reg[16]_0 ({core_n_1997,ptw_n_191,core_n_1998,core_n_1999}),
        .\reg_pmp_5_addr_reg[23] ({core_n_1935,core_n_1936,core_n_1937,core_n_1938}),
        .\reg_pmp_5_addr_reg[24] ({core_n_1911,core_n_1912,core_n_1913,core_n_1914}),
        .\reg_pmp_5_addr_reg[29] ({core_n_1850,core_n_1851,core_n_1852}),
        .\reg_pmp_5_addr_reg[4] (core_n_2033),
        .\reg_pmp_5_addr_reg[7] ({core_n_2025,core_n_2026,core_n_2027,core_n_2028}),
        .\reg_pmp_5_addr_reg[8] ({core_n_2029,core_n_2030,core_n_2031,core_n_2032}),
        .\reg_pmp_5_addr_reg[8]_0 ({frontend_io_ptw_pmp_5_addr[8:5],frontend_io_ptw_pmp_5_addr[3:0]}),
        .\reg_pmp_6_addr_reg[16] ({core_n_1975,core_n_1976,core_n_1977,core_n_1978}),
        .\reg_pmp_6_addr_reg[23] ({core_n_1928,core_n_1929,core_n_1930,core_n_1931}),
        .\reg_pmp_6_addr_reg[24] ({core_n_1919,core_n_1920,core_n_1921,core_n_1922}),
        .\reg_pmp_6_addr_reg[29] ({core_n_1844,core_n_1845,core_n_1846}),
        .\reg_pmp_6_addr_reg[2] (core_n_2069),
        .\reg_pmp_6_addr_reg[7] ({core_n_2061,core_n_2062,core_n_2063,core_n_2064}),
        .\reg_pmp_6_addr_reg[8] ({core_n_2065,core_n_2066,core_n_2067,core_n_2068}),
        .\reg_pmp_6_addr_reg[8]_0 ({frontend_io_ptw_pmp_6_addr[8:3],frontend_io_ptw_pmp_6_addr[1:0]}),
        .reg_pmp_6_cfg_w_reg(core_n_1836),
        .\reg_pmp_7_addr_reg[16] ({core_n_1971,core_n_1972,core_n_1973,core_n_1974}),
        .\reg_pmp_7_addr_reg[16]_0 ({core_n_1979,core_n_1980,core_n_1981,core_n_1982}),
        .\reg_pmp_7_addr_reg[23] ({core_n_1923,core_n_1924,core_n_1925,core_n_1926}),
        .\reg_pmp_7_addr_reg[24] ({core_n_1915,core_n_1916,core_n_1917,core_n_1918}),
        .\reg_pmp_7_addr_reg[29] ({core_n_1847,core_n_1848,core_n_1849}),
        .\reg_pmp_7_addr_reg[6] (core_n_2078),
        .\reg_pmp_7_addr_reg[7] ({core_n_2070,core_n_2071,core_n_2072,core_n_2073}),
        .\reg_pmp_7_addr_reg[8] ({core_n_2074,core_n_2075,core_n_2076,core_n_2077}),
        .\reg_pmp_7_addr_reg[8]_0 ({frontend_io_ptw_pmp_7_addr[8:7],frontend_io_ptw_pmp_7_addr[5:0]}),
        .\reg_sbadaddr_reg[30] (dcache_n_558),
        .\reg_scause_reg[1] (dcache_n_557),
        .release_ack_wait30_out(release_ack_wait30_out),
        .release_ack_wait_reg_0(dcache_n_90),
        .release_ack_wait_reg_1(sync_xing_n_207),
        .\remainder_reg[94] (div_io_resp_bits_data),
        .\req_tag_reg[4] (div_io_resp_bits_tag),
        .resp_ae_reg(ptw_n_132),
        .resp_ae_reg_0(core_n_649),
        .resp_valid_0_reg(ptw_n_193),
        .resp_valid_0_reg_0(ptw_n_195),
        .resp_valid_0_reg_1(ptw_n_196),
        .resp_valid_0_reg_2(ptw_n_197),
        .resp_valid_0_reg_3(ptw_n_131),
        .s0_clk_en(s0_clk_en),
        .s1_kill_reg(ptw_n_73),
        .s1_probe_reg_0(dcache_n_346),
        .s1_probe_reg_1(dcache_n_415),
        .s1_release_data_valid(s1_release_data_valid),
        .\s1_req_addr_reg[11]_0 (ptw_n_138),
        .\s1_req_addr_reg[11]_1 (ptw_n_145),
        .\s1_req_addr_reg[11]_2 (ptw_n_149),
        .\s1_req_addr_reg[11]_3 (ptw_n_156),
        .\s1_req_addr_reg[11]_4 (ptw_n_158),
        .\s1_req_addr_reg[2]_0 (ptw_n_152),
        .\s1_req_addr_reg[2]_1 (ptw_n_137),
        .\s1_req_addr_reg[2]_2 (ptw_n_148),
        .\s1_req_addr_reg[2]_3 (ptw_n_155),
        .\s1_req_addr_reg[32]_0 ({ptw_n_135,ptw_n_136}),
        .\s1_req_addr_reg[32]_1 ({ptw_n_164,ptw_n_165}),
        .\s1_req_addr_reg[39]_0 (dcache_n_416),
        .s1_req_phys_reg_0(core_n_423),
        .s1_req_phys_reg_1(\tlb/_T_194 ),
        .s1_req_phys_reg_2(\tlb/_T_210 ),
        .s1_valid(s1_valid),
        .s1_valid_reg_0(sync_xing_n_34),
        .\s2_data_reg[15]_0 ({dcache_n_17,dcache_n_18,dcache_n_19,dcache_n_20,dcache_n_21,dcache_n_22,dcache_n_23,dcache_n_24}),
        .\s2_data_reg[23]_0 ({dcache_n_25,dcache_n_26,dcache_n_27,dcache_n_28,dcache_n_29,dcache_n_30,dcache_n_31,dcache_n_32}),
        .\s2_data_reg[31]_0 ({dcache_n_33,dcache_n_34,dcache_n_35,dcache_n_36,dcache_n_37,dcache_n_38,dcache_n_39,dcache_n_40}),
        .\s2_data_reg[39]_0 ({dcache_n_41,dcache_n_42,dcache_n_43,dcache_n_44,dcache_n_45,dcache_n_46,dcache_n_47,dcache_n_48}),
        .\s2_data_reg[47]_0 ({dcache_n_49,dcache_n_50,dcache_n_51,dcache_n_52,dcache_n_53,dcache_n_54,dcache_n_55,dcache_n_56}),
        .\s2_data_reg[55]_0 ({dcache_n_57,dcache_n_58,dcache_n_59,dcache_n_60,dcache_n_61,dcache_n_62,dcache_n_63,dcache_n_64}),
        .\s2_data_reg[63]_0 ({dcache_n_65,dcache_n_66,dcache_n_67,dcache_n_68,dcache_n_69,dcache_n_70,dcache_n_71,dcache_n_72}),
        .\s2_data_reg[63]_1 (dcache_n_423),
        .s2_release_data_valid0(s2_release_data_valid0),
        .\s2_req_addr_reg[30]_0 (dcache_n_89),
        .s2_uncached(s2_uncached),
        .\size_reg[1] (tlMasterXbar_auto_out_a_bits_size[1]),
        .state(\tlb/state ),
        .state_0(\tlb/state_2 ),
        .\state_reg[0] (dcache_n_576),
        .\state_reg[0]_0 (dcache_n_578),
        .\state_reg[0]_1 (ptw_n_2),
        .\state_reg[0]_2 (ptw_n_52),
        .\state_reg[0]_3 (ptw_n_72),
        .\state_reg[1] (ptw_n_55),
        .\state_reg[1]_0 (ptw_n_1),
        .\state_reg[1]_1 (p_4_in),
        .\state_reg[1]_2 (ptw_n_16),
        .sys_reset_reg(sync_xing_n_350),
        .tag_array_0_reg_0(dcache_n_436),
        .target_reset(target_reset),
        .tlMasterXbar_auto_in_0_a_bits_size(tlMasterXbar_auto_in_0_a_bits_size),
        .tlMasterXbar_auto_in_0_d_bits_error(tlMasterXbar_auto_in_0_d_bits_error),
        .tlMasterXbar_auto_in_0_d_bits_size(tlMasterXbar_auto_in_0_d_bits_size),
        .tlMasterXbar_auto_out_b_bits_source(tlMasterXbar_auto_out_b_bits_source),
        .tlb_io_req_bits_sfence_bits_rs2(tlb_io_req_bits_sfence_bits_rs2),
        .traverse(traverse),
        .\uncachedReqs_0_addr_reg[2]_0 (dcache_n_210),
        .\uncachedReqs_0_tag_reg[6]_0 (dcacheArb_io_requestor_1_resp_bits_tag),
        .\valid_reg[0] (dcache_n_634),
        .\valid_reg[2] (core_n_1840),
        .\valid_reg[3] (dcache_n_429),
        .value(\Queue_3/value ),
        .value_1(\Queue_3/value_1 ),
        .value_1_reg(sync_xing_n_359),
        .value_1_reg_0(sync_xing_n_42),
        .value_1_reg_1(sync_xing_n_357),
        .value_1_reg_2(sync_xing_n_352),
        .value_1_reg_3(sync_xing_n_358),
        .value_1_reg_4(sync_xing_n_356),
        .value_1_reg_5(sync_xing_n_354),
        .value_1_reg_6(sync_xing_n_355),
        .value_1_reg_7(tlMasterXbar_auto_in_0_b_bits_size),
        .value_reg(sync_xing_n_220),
        .value_reg_0(sync_xing_n_209),
        .value_reg_1(sync_xing_n_208),
        .value_reg_2(sync_xing_n_50),
        .wb_ctrl_mem(wb_ctrl_mem),
        .wb_ctrl_mem_reg(core_n_1343),
        .\wb_reg_cause_reg[63] (core_n_1778),
        .\wb_reg_cause_reg[63]_0 (_T_2504),
        .\wb_reg_cause_reg[63]_1 (_T_2507),
        .\wb_reg_cause_reg[63]_2 (_T_2422),
        .\wb_reg_inst_reg[10] (wb_waddr[3]),
        .wb_reg_replay(wb_reg_replay),
        .wb_reg_valid(wb_reg_valid),
        .wb_reg_valid_reg(core_n_1344));
  HellaCacheArbiter dcacheArb
       (.Q(dcache_io_ptw_resp_bits_pte_ppn),
        ._T_177(_T_177),
        ._T_179(_T_179),
        .dcacheArb_io_requestor_0_req_bits_addr(dcacheArb_io_requestor_0_req_bits_addr),
        .dcacheArb_io_requestor_1_req_bits_addr(dcacheArb_io_requestor_1_req_bits_addr[31:3]),
        .dcache_io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),
        .host_clk(host_clk),
        .\state_reg[0] (ptw_n_2),
        .\state_reg[1] (p_4_in),
        .\state_reg[1]_0 (ptw_n_1));
  Frontend frontend
       (.ADDRA(_T_1396__T_1415_addr),
        .ADDRARDADDR({sync_xing_n_54,sync_xing_n_55,sync_xing_n_56,sync_xing_n_57,sync_xing_n_58,sync_xing_n_59}),
        .ADDRBWRADDR(ADDRBWRADDR[8:1]),
        .CO(\tlb/_T_384 ),
        .D(\tlb/_GEN_29 ),
        .DOA(tlMasterXbar_auto_in_0_d_bits_opcode),
        .E(sync_xing_n_41),
        .Q(tlMasterXbar_auto_in_1_a_bits_address),
        .S(frontend_n_92),
        .SR(\icache/p_0_in ),
        .WEBWE(sync_xing_n_40),
        ._GEN_274(_GEN_274[31:2]),
        ._GEN_55(_GEN_55),
        ._GEN_61(_GEN_61),
        ._T_100(\ibuf/_T_100 ),
        ._T_1005({_T_1005[6],_T_1005[4]}),
        ._T_1031({_T_1031[14],_T_1031[3]}),
        ._T_1050({_T_1050[5],_T_1050[2]}),
        ._T_1081(\tlb/_T_1081 ),
        ._T_1142({_T_1142[30],_T_1142[13:12]}),
        ._T_1406(_T_1406[31:2]),
        ._T_1573(_T_1573),
        ._T_1790(_T_1790),
        ._T_1821(_T_1821),
        .\_T_191_reg[0] (ADDRBWRADDR[0]),
        .\_T_191_reg[3] (\icache/_T_191_reg__0 ),
        .\_T_191_reg[6] (frontend_n_243),
        ._T_200__0({\tlb/_T_200__0 [30:29],\tlb/_T_200__0 [24:17],\tlb/_T_200__0 [15:14],\tlb/_T_200__0 [12]}),
        ._T_215_reg_0(core_n_686),
        .\_T_2547_reg[16] (_T_2549),
        .\_T_2547_reg[29] (core_n_1099),
        .\_T_2547_reg[31] (core_n_1100),
        ._T_382(\tlb/_T_382 ),
        ._T_382__0({\tlb/_T_382__0 [28:27],\tlb/_T_382__0 [25]}),
        ._T_480(\tlb/_T_480 ),
        ._T_726(\tlb/_T_726 ),
        ._T_877(_T_877),
        ._T_889({_T_889[24:15],_T_889[11:7]}),
        ._T_909({_T_909[31],_T_909[29:26]}),
        .\_T_973_reg[2] (\tlb/_T_1432 ),
        .bad_va(\tlb/bad_va ),
        .\buf__data_reg[0] (core__86_n_0),
        .\buf__data_reg[0]_0 (core__71_n_0),
        .\buf__data_reg[0]_1 (core__85_n_0),
        .\buf__data_reg[10] (core__69_n_0),
        .\buf__data_reg[12] (core__53_n_0),
        .\buf__data_reg[12]_0 (core__50_n_0),
        .\buf__data_reg[12]_1 (core__52_n_0),
        .\buf__data_reg[12]_2 (core__58_n_0),
        .\buf__data_reg[12]_3 (core__45_n_0),
        .\buf__data_reg[12]_4 (core__40_n_0),
        .\buf__data_reg[12]_5 (core__59_n_0),
        .\buf__data_reg[13] (core__60_n_0),
        .\buf__data_reg[13]_0 (core__76_n_0),
        .\buf__data_reg[14] ({frontend_io_cpu_resp_bits_data[30:28],frontend_io_cpu_resp_bits_data[26],frontend_io_cpu_resp_bits_data[23],frontend_io_cpu_resp_bits_data[19],frontend_io_cpu_resp_bits_data[14:12],frontend_io_cpu_resp_bits_data[10],frontend_io_cpu_resp_bits_data[7],frontend_io_cpu_resp_bits_data[3]}),
        .\buf__data_reg[14]_0 (core__66_n_0),
        .\buf__data_reg[14]_1 (core__84_n_0),
        .\buf__data_reg[14]_2 (core__78_n_0),
        .\buf__data_reg[14]_3 (core__57_n_0),
        .\buf__data_reg[14]_4 (core__79_n_0),
        .\buf__data_reg[15] (\ibuf/_T_74 ),
        .\buf__data_reg[15]_0 (core__70_n_0),
        .\buf__data_reg[15]_1 (core__68_n_0),
        .\buf__data_reg[15]_2 (core__88_n_0),
        .\buf__data_reg[15]_3 (core__75_n_0),
        .\buf__data_reg[15]_4 (core__89_n_0),
        .\buf__data_reg[15]_5 ({core_n_2086,core_n_2087,core_n_2088,core_n_2089,core_n_2090,core_n_2091,core_n_2092,core_n_2093,core_n_2094,core_n_2095,core_n_2096,core_n_2097,core_n_2098,core_n_2099,core_n_2100,core_n_2101}),
        .\buf__data_reg[15]_6 (core__72_n_0),
        .\buf__data_reg[15]_7 (core_n_1238),
        .\buf__data_reg[1] (core__61_n_0),
        .\buf__data_reg[1]_0 (core__90_n_0),
        .\buf__data_reg[1]_1 (core__65_n_0),
        .\buf__data_reg[1]_10 (core__51_n_0),
        .\buf__data_reg[1]_2 (core__83_n_0),
        .\buf__data_reg[1]_3 (core__82_n_0),
        .\buf__data_reg[1]_4 (core__46_n_0),
        .\buf__data_reg[1]_5 (core__697_n_0),
        .\buf__data_reg[1]_6 (core__56_n_0),
        .\buf__data_reg[1]_7 (core__699_n_0),
        .\buf__data_reg[1]_8 (core_n_1098),
        .\buf__data_reg[1]_9 (core__702_n_0),
        .\buf__data_reg[2] (core__54_n_0),
        .\buf__data_reg[3] (core__81_n_0),
        .\buf__data_reg[3]_0 (core__62_n_0),
        .\buf__data_reg[3]_1 (core__714_n_0),
        .\buf__data_reg[3]_2 (core__39_n_0),
        .\buf__data_reg[3]_3 (core__695_n_0),
        .\buf__data_reg[3]_4 (core__41_n_0),
        .\buf__data_reg[4] (core__64_n_0),
        .\buf__data_reg[4]_0 (core__43_n_0),
        .\buf__data_reg[5] (core__74_n_0),
        .\buf__data_reg[6] (core__80_n_0),
        .\buf__data_reg[7] (core__42_n_0),
        .\buf__data_reg[9] (core__63_n_0),
        .buf__pc(\ibuf/buf__pc ),
        .\buf__pc_reg[1] (frontend_n_265),
        .\buf__pc_reg[1]_0 (\ibuf/_T_81 ),
        .\buf__pc_reg[39] ({core_n_1069,core_n_1070,core_n_1071,core_n_1072,core_n_1073,core_n_1074,core_n_1075,core_n_1076,core_n_1077,core_n_1078,core_n_1079,core_n_1080,core_n_1081,core_n_1082,core_n_1083,core_n_1084,core_n_1085,core_n_1086,core_n_1087}),
        .buf__replay(\ibuf/buf__replay ),
        .buf__xcpt_ae_inst(\ibuf/buf__xcpt_ae_inst ),
        .buf__xcpt_pf_inst_reg(core_n_1256),
        .buf__xcpt_pf_inst_reg_0(core_n_95),
        .data_arrays_0_0_reg(frontend_n_240),
        .data_arrays_0_0_reg_0(frontend_n_241),
        .data_arrays_0_0_reg_i_20__0(data_arrays_0_0_reg_i_20__0),
        .data_arrays_0_0_reg_i_21__0(data_arrays_0_0_reg_i_21__0),
        .data_arrays_0_0_reg_i_22__0(data_arrays_0_0_reg_i_22__0),
        .data_arrays_0_0_reg_i_23__0(data_arrays_0_0_reg_i_23__0),
        .data_arrays_0_0_reg_i_24__0(data_arrays_0_0_reg_i_24__0),
        .data_arrays_0_0_reg_i_25__0(data_arrays_0_0_reg_i_25__0),
        .data_arrays_0_0_reg_i_26__0(data_arrays_0_0_reg_i_26__0),
        .data_arrays_0_0_reg_i_27__0(data_arrays_0_0_reg_i_27__0),
        .data_arrays_0_0_reg_i_28__0(data_arrays_0_0_reg_i_28__0),
        .data_arrays_1_0_reg_i_11(data_arrays_1_0_reg_i_11),
        .data_arrays_1_0_reg_i_12(data_arrays_1_0_reg_i_12),
        .data_arrays_1_0_reg_i_13(data_arrays_1_0_reg_i_13),
        .data_arrays_1_0_reg_i_14(data_arrays_1_0_reg_i_14),
        .data_arrays_1_0_reg_i_15(data_arrays_1_0_reg_i_15),
        .data_arrays_1_0_reg_i_16(data_arrays_1_0_reg_i_16),
        .data_arrays_1_0_reg_i_17(data_arrays_1_0_reg_i_17),
        .data_arrays_1_0_reg_i_18(data_arrays_1_0_reg_i_18),
        .data_arrays_1_0_reg_i_19(data_arrays_1_0_reg_i_19),
        .dcache_blocked_reg(core_n_1090),
        .dcache_io_ptw_resp_bits_level(dcache_io_ptw_resp_bits_level),
        .doUncachedResp_reg(core_n_1092),
        .\elts_4_pc_reg[38] ({s2_pc[38],s2_pc[1]}),
        .\ex_ctrl_alu_fn_reg[3] (id_ctrl_alu_fn),
        .\ex_ctrl_csr_reg[0] (frontend_n_225),
        .\ex_ctrl_csr_reg[1] (frontend_n_231),
        .\ex_ctrl_csr_reg[1]_0 ({core_n_92,core_n_93}),
        .ex_ctrl_div_reg(frontend_n_404),
        .ex_ctrl_fence_i_reg(frontend_n_396),
        .\ex_ctrl_mem_cmd_reg[2] (frontend_n_366),
        .\ex_ctrl_mem_cmd_reg[2]_0 (id_ctrl_mem_cmd[2:0]),
        .\ex_ctrl_mem_cmd_reg[2]_1 (frontend_n_386),
        .\ex_ctrl_mem_cmd_reg[4] (frontend_n_304),
        .ex_ctrl_mem_reg(frontend_n_318),
        .ex_ctrl_mem_reg_0(frontend_n_358),
        .ex_ctrl_mem_reg_1(frontend_n_365),
        .ex_ctrl_mem_reg_2(frontend_n_368),
        .ex_ctrl_mem_reg_3(frontend_n_369),
        .ex_ctrl_mem_reg_4(frontend_n_370),
        .ex_ctrl_mem_reg_5(frontend_n_387),
        .ex_ctrl_mem_reg_6(frontend_n_391),
        .ex_ctrl_mem_reg_7(frontend_n_403),
        .\ex_ctrl_mem_type_reg[0] (frontend_n_232),
        .\ex_ctrl_mem_type_reg[1] ({frontend_n_359,frontend_n_360}),
        .\ex_ctrl_mem_type_reg[1]_0 (frontend_n_361),
        .\ex_ctrl_mem_type_reg[1]_1 (frontend_n_362),
        .\ex_ctrl_mem_type_reg[1]_2 (frontend_n_371),
        .ex_ctrl_rxs2_reg(frontend_n_367),
        .\ex_ctrl_sel_alu1_reg[0] (frontend_n_390),
        .\ex_ctrl_sel_alu2_reg[0] (frontend_n_356),
        .\ex_ctrl_sel_alu2_reg[0]_0 (frontend_n_392),
        .\ex_ctrl_sel_alu2_reg[0]_1 (frontend_n_419),
        .\ex_ctrl_sel_alu2_reg[1] (frontend_n_169),
        .\ex_ctrl_sel_alu2_reg[1]_0 (frontend_n_170),
        .\ex_ctrl_sel_alu2_reg[1]_1 (frontend_n_222),
        .\ex_ctrl_sel_alu2_reg[1]_10 (frontend_n_395),
        .\ex_ctrl_sel_alu2_reg[1]_11 (frontend_n_402),
        .\ex_ctrl_sel_alu2_reg[1]_12 (frontend_n_409),
        .\ex_ctrl_sel_alu2_reg[1]_2 (frontend_n_223),
        .\ex_ctrl_sel_alu2_reg[1]_3 (frontend_n_224),
        .\ex_ctrl_sel_alu2_reg[1]_4 (frontend_n_352),
        .\ex_ctrl_sel_alu2_reg[1]_5 (frontend_n_354),
        .\ex_ctrl_sel_alu2_reg[1]_6 (frontend_n_355),
        .\ex_ctrl_sel_alu2_reg[1]_7 (frontend_n_378),
        .\ex_ctrl_sel_alu2_reg[1]_8 (frontend_n_389),
        .\ex_ctrl_sel_alu2_reg[1]_9 (frontend_n_393),
        .\ex_ctrl_sel_imm_reg[2] (frontend_n_312),
        .\ex_ctrl_sel_imm_reg[2]_0 (id_ctrl_sel_imm[2]),
        .ex_ctrl_wxd_reg(frontend_n_364),
        .ex_ctrl_wxd_reg_0(core_n_1102),
        .ex_ctrl_wxd_reg_1(core_n_1362),
        .ex_reg_flush_pipe_reg(frontend_n_226),
        .ex_reg_flush_pipe_reg_0(frontend_n_230),
        .\ex_reg_inst_reg[10] (frontend_n_268),
        .\ex_reg_inst_reg[10]_0 (frontend_n_269),
        .\ex_reg_inst_reg[10]_1 (core_n_1240),
        .\ex_reg_inst_reg[11] (dcacheArb_io_requestor_1_req_bits_tag),
        .\ex_reg_inst_reg[14] (frontend_n_293),
        .\ex_reg_inst_reg[23] (frontend_n_300),
        .\ex_reg_inst_reg[24] (frontend_n_285),
        .\ex_reg_inst_reg[24]_0 (frontend_n_294),
        .\ex_reg_inst_reg[29] ({ibuf_io_inst_0_bits_raw[29],ibuf_io_inst_0_bits_raw[25],ibuf_io_inst_0_bits_raw[22],ibuf_io_inst_0_bits_raw[15:14],ibuf_io_inst_0_bits_raw[12:11],ibuf_io_inst_0_bits_raw[9:8],ibuf_io_inst_0_bits_raw[6:0]}),
        .\ex_reg_inst_reg[31] (frontend_n_267),
        .ex_reg_load_use_reg(frontend_n_372),
        .ex_reg_load_use_reg_0(frontend_n_374),
        .ex_reg_load_use_reg_1(frontend_n_376),
        .ex_reg_load_use_reg_2(frontend_n_410),
        .\ex_reg_pc_reg[38] (\fq/elts_0_pc ),
        .\ex_reg_pc_reg[39] ({ibuf_io_pc[39:37],ibuf_io_pc[35],ibuf_io_pc[33],ibuf_io_pc[31],ibuf_io_pc[29],ibuf_io_pc[27],ibuf_io_pc[25],ibuf_io_pc[23],ibuf_io_pc[21],ibuf_io_pc[19],ibuf_io_pc[17],ibuf_io_pc[15],ibuf_io_pc[13],ibuf_io_pc[11],ibuf_io_pc[9],ibuf_io_pc[7],ibuf_io_pc[5]}),
        .\ex_reg_pc_reg[5] (frontend_n_54),
        .ex_reg_rs_bypass_1_reg(frontend_n_375),
        .\ex_reg_rs_lsb_0_reg[0] (frontend_n_353),
        .\ex_reg_rs_lsb_0_reg[0]_0 (frontend_n_373),
        .\ex_reg_rs_msb_0_reg[29] (p_1_in),
        .\ex_reg_rs_msb_0_reg[29]_0 (frontend_n_351),
        .\ex_reg_rs_msb_0_reg[59] (_T_1396__T_1405_addr),
        .\ex_reg_rs_msb_0_reg[61] (frontend_n_388),
        .\ex_reg_rs_msb_1_reg[61] (frontend_n_416),
        .fq_reset(fq_reset),
        .frontend_io_cpu_req_bits_speculative(frontend_io_cpu_req_bits_speculative),
        .frontend_io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
        .frontend_io_cpu_resp_bits_replay(frontend_io_cpu_resp_bits_replay),
        .frontend_io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),
        .frontend_io_cpu_resp_bits_xcpt_pf_inst(frontend_io_cpu_resp_bits_xcpt_pf_inst),
        .frontend_io_cpu_resp_valid(frontend_io_cpu_resp_valid),
        .frontend_io_cpu_sfence_valid(frontend_io_cpu_sfence_valid),
        .frontend_io_ptw_ptbr_mode(frontend_io_ptw_ptbr_mode),
        .frontend_io_ptw_req_ready(frontend_io_ptw_req_ready),
        .frontend_io_ptw_status_prv(frontend_io_ptw_status_prv),
        .hitsVec_4(\tlb/hitsVec_4 ),
        .host_clk(host_clk),
        .ibuf_io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
        .ibuf_io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
        .ibuf_io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
        .id_ctrl_alu_dw(id_ctrl_alu_dw),
        .id_ctrl_fence_i(id_ctrl_fence_i),
        .id_ctrl_jal(id_ctrl_jal),
        .id_ctrl_mem(id_ctrl_mem),
        .id_ctrl_rxs2(id_ctrl_rxs2),
        .id_ctrl_sel_alu1(id_ctrl_sel_alu1[1]),
        .id_ctrl_wxd(id_ctrl_wxd),
        .id_reg_fence_reg(core_n_1091),
        .invalidated(\icache/invalidated ),
        .invalidated_reg(sync_xing_n_35),
        .invalidated_reg_0(sync_xing_n_39),
        .io_mask(fq_io_mask),
        .lastGrant(\arb/lastGrant ),
        .load(\icache/load ),
        .mem_ctrl_mem(mem_ctrl_mem),
        .\mem_reg_inst_reg[11] ({mem_waddr[4],mem_waddr[2]}),
        .\mem_reg_inst_reg[9] (core_n_1094),
        .mem_reg_valid_reg(mem_reg_replay_reg),
        .nBufValid_reg(frontend_n_320),
        .nBufValid_reg_0(core__97_n_0),
        .nBufValid_reg_1(core__99_n_0),
        .nBufValid_reg_10(core__93_n_0),
        .nBufValid_reg_11(core__47_n_0),
        .nBufValid_reg_12(core__698_n_0),
        .nBufValid_reg_2(core__98_n_0),
        .nBufValid_reg_3(core_n_892),
        .nBufValid_reg_4(core__73_n_0),
        .nBufValid_reg_5(core__67_n_0),
        .nBufValid_reg_6(core__91_n_0),
        .nBufValid_reg_7(core__92_n_0),
        .nBufValid_reg_8(core__87_n_0),
        .nBufValid_reg_9(core__77_n_0),
        .p_12_in(\icache/p_12_in ),
        .p_13_in(\tlb/p_13_in ),
        .p_2_in(\tlb/p_2_in ),
        .p_31_in(p_31_in),
        .\r_pte_ppn_reg[16] (ptw_n_53),
        .\r_pte_ppn_reg[19] (dcache_io_ptw_resp_bits_pte_ppn),
        .r_pte_u_reg({dcache_io_ptw_resp_bits_pte_u,dcache_io_ptw_resp_bits_pte_g,dcache_io_ptw_resp_bits_ae,\tlb/_T_943_4 ,\tlb/_T_952 }),
        .\r_refill_tag_reg[26] (dcache_io_ptw_req_bits_addr),
        .\r_refill_waddr_reg[1] (\tlb/_T_815 ),
        .\r_refill_waddr_reg[1]_0 (core_n_685),
        .\r_req_addr_reg[26] (arb_io_out_bits_addr),
        .r_req_dest_reg(frontend_n_44),
        .ram_data__T_63_data(tlMasterXbar_auto_in_0_d_bits_data),
        .refill_one_beat(\icache/refill_one_beat ),
        .refill_valid(\icache/refill_valid ),
        .refill_valid_reg(frontend_n_49),
        .\reg_bp_0_address_reg[38] (csr_io_bp_0_address[38]),
        .\reg_bp_0_control_tmatch_reg[1] (core_n_1089),
        .reg_debug_reg(core_n_890),
        .\reg_entries_0_reg[0] ({\tlb/p_0_in_1 [19],\tlb/p_0_in_1 [16],\tlb/p_0_in_1 [13]}),
        .\reg_entries_0_reg[0]_0 (frontend_n_126),
        .\reg_entries_0_reg[5] (\tlb/pmp/_T_53 ),
        .\reg_entries_0_reg[5]_0 (\tlb/pmp/_T_58 ),
        .\reg_entries_0_reg[5]_1 (\tlb/pmp/_T_89 ),
        .\reg_entries_0_reg[5]_10 (frontend_n_117),
        .\reg_entries_0_reg[5]_11 (frontend_n_118),
        .\reg_entries_0_reg[5]_12 (frontend_n_119),
        .\reg_entries_0_reg[5]_13 (frontend_n_120),
        .\reg_entries_0_reg[5]_14 (frontend_n_121),
        .\reg_entries_0_reg[5]_15 (frontend_n_125),
        .\reg_entries_0_reg[5]_16 (frontend_n_127),
        .\reg_entries_0_reg[5]_17 (frontend_n_128),
        .\reg_entries_0_reg[5]_18 (frontend_n_129),
        .\reg_entries_0_reg[5]_19 (frontend_n_130),
        .\reg_entries_0_reg[5]_2 (\tlb/pmp/_T_125 ),
        .\reg_entries_0_reg[5]_20 (frontend_n_131),
        .\reg_entries_0_reg[5]_21 (frontend_n_132),
        .\reg_entries_0_reg[5]_22 (frontend_n_133),
        .\reg_entries_0_reg[5]_23 (frontend_n_134),
        .\reg_entries_0_reg[5]_24 (frontend_n_136),
        .\reg_entries_0_reg[5]_25 (frontend_n_137),
        .\reg_entries_0_reg[5]_26 (frontend_n_138),
        .\reg_entries_0_reg[5]_27 (frontend_n_139),
        .\reg_entries_0_reg[5]_28 (frontend_n_140),
        .\reg_entries_0_reg[5]_29 (frontend_n_141),
        .\reg_entries_0_reg[5]_3 (\tlb/pmp/_T_161 ),
        .\reg_entries_0_reg[5]_30 (frontend_n_142),
        .\reg_entries_0_reg[5]_31 (frontend_n_143),
        .\reg_entries_0_reg[5]_32 (frontend_n_144),
        .\reg_entries_0_reg[5]_33 (frontend_n_145),
        .\reg_entries_0_reg[5]_34 (frontend_n_146),
        .\reg_entries_0_reg[5]_35 (frontend_n_147),
        .\reg_entries_0_reg[5]_36 (frontend_n_148),
        .\reg_entries_0_reg[5]_37 (frontend_n_149),
        .\reg_entries_0_reg[5]_38 (frontend_n_150),
        .\reg_entries_0_reg[5]_39 (frontend_n_151),
        .\reg_entries_0_reg[5]_4 (\tlb/pmp/_T_197 ),
        .\reg_entries_0_reg[5]_40 (frontend_n_152),
        .\reg_entries_0_reg[5]_5 (\tlb/pmp/_T_233 ),
        .\reg_entries_0_reg[5]_6 (\tlb/pmp/_T_269 ),
        .\reg_entries_0_reg[5]_7 (frontend_n_114),
        .\reg_entries_0_reg[5]_8 (frontend_n_115),
        .\reg_entries_0_reg[5]_9 (frontend_n_116),
        .\reg_entries_1_reg[0] ({frontend_n_51,frontend_n_52}),
        .\reg_misa_reg[12] (csr_io_status_isa[12]),
        .\reg_misa_reg[2] (core_n_1097),
        .\reg_mstatus_prv_reg[1] (core_n_752),
        .reg_mstatus_tsr_reg(core_n_70),
        .reg_mstatus_tvm_reg(core__94_n_0),
        .reg_mstatus_tw_reg(core_n_69),
        .\reg_pmp_0_addr_reg[14] ({core_n_745,core_n_746,core_n_747,core_n_748}),
        .\reg_pmp_0_addr_reg[22] ({core_n_805,core_n_806,core_n_807,core_n_808}),
        .\reg_pmp_0_addr_reg[28] ({core_n_753,core_n_754,core_n_755}),
        .\reg_pmp_0_addr_reg[29] (frontend_io_ptw_pmp_0_addr[29:10]),
        .\reg_pmp_0_addr_reg[6] ({core_n_815,core_n_816,core_n_817,core_n_818}),
        .\reg_pmp_0_addr_reg[6]_0 ({core_n_811,core_n_812,core_n_813,core_n_814}),
        .\reg_pmp_0_addr_reg[8] (core_n_819),
        .\reg_pmp_1_addr_reg[14] ({core_n_736,core_n_737,core_n_738,core_n_739}),
        .\reg_pmp_1_addr_reg[22] ({core_n_801,core_n_802,core_n_803,core_n_804}),
        .\reg_pmp_1_addr_reg[28] ({core_n_756,core_n_757,core_n_758}),
        .\reg_pmp_1_addr_reg[29] (frontend_io_ptw_pmp_1_addr[29:10]),
        .\reg_pmp_1_addr_reg[6] ({core_n_824,core_n_825,core_n_826,core_n_827}),
        .\reg_pmp_1_addr_reg[6]_0 ({core_n_820,core_n_821,core_n_822,core_n_823}),
        .\reg_pmp_1_addr_reg[8] (core_n_828),
        .\reg_pmp_2_addr_reg[14] ({core_n_730,core_n_731,core_n_732,core_n_733}),
        .\reg_pmp_2_addr_reg[22] ({core_n_797,core_n_798,core_n_799,core_n_800}),
        .\reg_pmp_2_addr_reg[28] ({core_n_759,core_n_760,core_n_761}),
        .\reg_pmp_2_addr_reg[29] (frontend_io_ptw_pmp_2_addr[29:10]),
        .\reg_pmp_2_addr_reg[6] ({core_n_833,core_n_834,core_n_835,core_n_836}),
        .\reg_pmp_2_addr_reg[6]_0 ({core_n_829,core_n_830,core_n_831,core_n_832}),
        .\reg_pmp_2_addr_reg[8] (core_n_837),
        .\reg_pmp_3_addr_reg[14] ({core_n_708,core_n_709,core_n_710,core_n_711}),
        .\reg_pmp_3_addr_reg[22] ({core_n_785,core_n_786,core_n_787,core_n_788}),
        .\reg_pmp_3_addr_reg[28] ({core_n_768,core_n_769,core_n_770}),
        .\reg_pmp_3_addr_reg[29] (frontend_io_ptw_pmp_3_addr[29:10]),
        .\reg_pmp_3_addr_reg[6] ({core_n_860,core_n_861,core_n_862,core_n_863}),
        .\reg_pmp_3_addr_reg[6]_0 ({core_n_856,core_n_857,core_n_858,core_n_859}),
        .\reg_pmp_3_addr_reg[8] (core_n_864),
        .\reg_pmp_4_addr_reg[14] ({core_n_700,core_n_701,core_n_702,core_n_703}),
        .\reg_pmp_4_addr_reg[22] ({core_n_781,core_n_782,core_n_783,core_n_784}),
        .\reg_pmp_4_addr_reg[28] ({core_n_771,core_n_772,core_n_773}),
        .\reg_pmp_4_addr_reg[29] (frontend_io_ptw_pmp_4_addr[29:10]),
        .\reg_pmp_4_addr_reg[6] ({core_n_869,core_n_870,core_n_871,core_n_872}),
        .\reg_pmp_4_addr_reg[6]_0 ({core_n_865,core_n_866,core_n_867,core_n_868}),
        .\reg_pmp_4_addr_reg[8] (core_n_873),
        .\reg_pmp_5_addr_reg[14] ({core_n_692,core_n_693,core_n_694,core_n_695}),
        .\reg_pmp_5_addr_reg[22] ({core_n_777,core_n_778,core_n_779,core_n_780}),
        .\reg_pmp_5_addr_reg[28] ({core_n_774,core_n_775,core_n_776}),
        .\reg_pmp_5_addr_reg[29] (frontend_io_ptw_pmp_5_addr[29:10]),
        .\reg_pmp_5_addr_reg[6] ({core_n_878,core_n_879,core_n_880,core_n_881}),
        .\reg_pmp_5_addr_reg[6]_0 ({core_n_874,core_n_875,core_n_876,core_n_877}),
        .\reg_pmp_5_addr_reg[8] (core_n_882),
        .\reg_pmp_6_addr_reg[14] ({core_n_721,core_n_722,core_n_723,core_n_724}),
        .\reg_pmp_6_addr_reg[22] ({core_n_793,core_n_794,core_n_795,core_n_796}),
        .\reg_pmp_6_addr_reg[28] ({core_n_762,core_n_763,core_n_764}),
        .\reg_pmp_6_addr_reg[29] (frontend_io_ptw_pmp_6_addr[29:10]),
        .\reg_pmp_6_addr_reg[6] ({core_n_842,core_n_843,core_n_844,core_n_845}),
        .\reg_pmp_6_addr_reg[6]_0 ({core_n_838,core_n_839,core_n_840,core_n_841}),
        .\reg_pmp_6_addr_reg[8] (core_n_846),
        .\reg_pmp_7_addr_reg[14] ({core_n_712,core_n_713,core_n_714,core_n_715}),
        .\reg_pmp_7_addr_reg[22] ({core_n_789,core_n_790,core_n_791,core_n_792}),
        .\reg_pmp_7_addr_reg[28] ({core_n_765,core_n_766,core_n_767}),
        .\reg_pmp_7_addr_reg[29] (frontend_io_ptw_pmp_7_addr[29:10]),
        .\reg_pmp_7_addr_reg[6] ({core_n_851,core_n_852,core_n_853,core_n_854}),
        .\reg_pmp_7_addr_reg[6]_0 ({core_n_847,core_n_848,core_n_849,core_n_850}),
        .\reg_pmp_7_addr_reg[8] (core_n_855),
        .\req_tag_reg[4] (dcache_n_544),
        .\req_tag_reg[4]_0 (core_n_1323),
        .resp_ae_reg(core_n_687),
        .resp_ae_reg_0(core_n_649),
        .resp_valid_1_reg(s2_valid_reg),
        .resp_valid_1_reg_0(core_n_883),
        .resp_valid_1_reg_1(core_n_884),
        .resp_valid_1_reg_2(core_n_885),
        .resp_valid_1_reg_3(core_n_886),
        .resp_valid_1_reg_4(core_n_887),
        .resp_valid_1_reg_5(core_n_888),
        .resp_valid_1_reg_6(core_n_889),
        .resp_valid_1_reg_7(core_n_809),
        .\s1_pc_reg[11]_0 ({D,frontend_n_239}),
        .\s1_pc_reg[38]_0 (core_n_749),
        .\s2_pc_reg[1]_0 (core_n_1029),
        .\s2_pc_reg[39]_0 ({s1_pc[39:38],s1_pc[31],s1_pc[28],s1_pc[25],s1_pc[11:2]}),
        .s2_replay(s2_replay),
        .\s2_req_tag_reg[4] (core__48_n_0),
        .\s2_req_tag_reg[5] (dcache_n_543),
        .\s2_req_tag_reg[5]_0 (dcache_n_554),
        .state(\tlb/state_2 ),
        .state_0(\tlb/state ),
        .sys_reset_reg(core_n_682),
        .sys_reset_reg_0(sys_reset_reg),
        .tag_array_0_reg(frontend_n_244),
        .tag_array_0_reg_0(frontend_n_245),
        .target_reset(target_reset),
        .tlMasterXbar_auto_in_0_d_bits_error(tlMasterXbar_auto_in_0_d_bits_error),
        .tlMasterXbar_auto_in_0_d_bits_size(tlMasterXbar_auto_in_0_d_bits_size[3]),
        .valid_2_reg(core_n_647),
        .\valid_reg[3] (\tlb/entries_3_g ),
        .value_1_reg(sync_xing_n_43),
        .value_1_reg_0(sync_xing_n_42),
        .value_1_reg_1(sync_xing_n_44),
        .value_1_reg_2(sync_xing_n_46),
        .value_1_reg_3(sync_xing_n_45),
        .value_1_reg_4(sync_xing_n_47),
        .value_1_reg_5(sync_xing_n_48),
        .value_1_reg_6({\icache/p_0_in__0 [8],\icache/p_0_in__0 [6],\icache/p_0_in__0 [4],\icache/p_0_in__0 [0]}),
        .value_reg(sync_xing_n_33),
        .wb_ctrl_fence_i_reg(core_n_680),
        .\wb_ctrl_mem_type_reg[0] (frontend_io_cpu_sfence_bits_rs1),
        .wb_ctrl_wxd_reg(core_n_1360),
        .\wb_reg_inst_reg[10] (core_n_1128),
        .\wb_reg_inst_reg[10]_0 (core_n_1239),
        .\wb_reg_inst_reg[11] (core__44_n_0),
        .\wb_reg_inst_reg[11]_0 (wb_waddr),
        .\wb_reg_inst_reg[9] (_T_1396__T_2475_addr),
        .\wb_reg_pc_reg[39] (frontend_io_cpu_req_bits_pc),
        .wb_reg_valid_reg(core_n_551));
  CARRY4 mem_br_taken__reg_i_3
       (.CI(mem_br_taken__reg_i_4_n_0),
        .CO({\alu/_T_31 ,mem_br_taken__reg_i_3_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,core_n_2317,core__182_n_0}));
  CARRY4 mem_br_taken__reg_i_4
       (.CI(mem_br_taken__reg_i_6_n_0),
        .CO({mem_br_taken__reg_i_4_n_0,mem_br_taken__reg_i_4_n_1,mem_br_taken__reg_i_4_n_2,mem_br_taken__reg_i_4_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core__181_n_0,core__180_n_0,core__179_n_0,core__178_n_0}));
  CARRY4 mem_br_taken__reg_i_6
       (.CI(mem_br_taken__reg_i_7_n_0),
        .CO({mem_br_taken__reg_i_6_n_0,mem_br_taken__reg_i_6_n_1,mem_br_taken__reg_i_6_n_2,mem_br_taken__reg_i_6_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core__177_n_0,core__176_n_0,core__175_n_0,core__174_n_0}));
  CARRY4 mem_br_taken__reg_i_7
       (.CI(mem_br_taken__reg_i_8_n_0),
        .CO({mem_br_taken__reg_i_7_n_0,mem_br_taken__reg_i_7_n_1,mem_br_taken__reg_i_7_n_2,mem_br_taken__reg_i_7_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core__173_n_0,core__172_n_0,core__171_n_0,core__170_n_0}));
  CARRY4 mem_br_taken__reg_i_8
       (.CI(mem_br_taken__reg_i_9_n_0),
        .CO({mem_br_taken__reg_i_8_n_0,mem_br_taken__reg_i_8_n_1,mem_br_taken__reg_i_8_n_2,mem_br_taken__reg_i_8_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core__169_n_0,core__168_n_0,core__167_n_0,core__166_n_0}));
  CARRY4 mem_br_taken__reg_i_9
       (.CI(\<const0> ),
        .CO({mem_br_taken__reg_i_9_n_0,mem_br_taken__reg_i_9_n_1,mem_br_taken__reg_i_9_n_2,mem_br_taken__reg_i_9_n_3}),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core__165_n_0,core__164_n_0,core__163_n_0,core__162_n_0}));
  PTW ptw
       (.CO(_T_2774),
        .D({_T_273,ptw_n_49,ptw_n_50,ptw_n_51}),
        .E(_T_439),
        .O(alu_io_adder_out),
        .Q(dcache_io_ptw_resp_bits_pte_ppn),
        .S(ptw_n_190),
        .SR(core_n_1799),
        ._T_1156(_T_1156),
        ._T_1498(_T_1498),
        ._T_1701(_T_1701[8]),
        ._T_177(_T_177),
        ._T_177_reg(p_4_in),
        ._T_179_reg(dcache_n_578),
        .\_T_1883_reg[1] (dcache_io_ptw_status_dprv[1]),
        ._T_255(_T_255),
        ._T_384(_T_384),
        .\_T_407_0_reg[19]_0 (ptw_n_82),
        ._T_407_1(_T_407_1),
        ._T_407_4(_T_407_4),
        ._T_407_6(_T_407_6),
        .\_T_407_7_reg[0]_0 (ptw_n_76),
        .\_T_407_7_reg[19]_0 (ptw_n_83),
        ._T_435(_T_435),
        ._T_499(_T_499),
        ._T_931(_T_931),
        .\bypass_mux_2_reg[63] (_T_2772),
        .dataArb_io_in_2_valid(dataArb_io_in_2_valid),
        .data_arrays_0_0_reg(ptw_n_56),
        .data_arrays_0_0_reg_0(ptw_n_66),
        .data_arrays_0_0_reg_1(ptw_n_67),
        .data_arrays_0_0_reg_2(ptw_n_68),
        .data_arrays_0_0_reg_3(ptw_n_69),
        .data_arrays_0_0_reg_4(ptw_n_70),
        .dcacheArb_io_requestor_0_req_bits_addr(dcacheArb_io_requestor_0_req_bits_addr),
        .dcacheArb_io_requestor_0_req_ready(dcacheArb_io_requestor_0_req_ready),
        .dcacheArb_io_requestor_0_s1_kill(dcacheArb_io_requestor_0_s1_kill),
        .dcacheArb_io_requestor_1_req_bits_addr({dcacheArb_io_requestor_1_req_bits_addr[38:32],dcacheArb_io_requestor_1_req_bits_addr[11:6],dcacheArb_io_requestor_1_req_bits_addr[2:0]}),
        .dcacheArb_io_requestor_1_req_ready(dcacheArb_io_requestor_1_req_ready),
        .dcacheArb_io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),
        .dcacheArb_io_requestor_1_resp_bits_data(dcacheArb_io_requestor_1_resp_bits_data[7]),
        .dcacheArb_io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),
        .dcacheArb_io_requestor_1_s2_xcpt_ae_ld(dcacheArb_io_requestor_1_s2_xcpt_ae_ld),
        .dcache_io_ptw_resp_bits_homogeneous(dcache_io_ptw_resp_bits_homogeneous),
        .dcache_io_ptw_resp_bits_level(dcache_io_ptw_resp_bits_level),
        .dcache_io_ptw_resp_bits_pte_v(dcache_io_ptw_resp_bits_pte_v),
        .dcache_io_ptw_resp_valid(dcache_io_ptw_resp_valid),
        .doUncachedResp_reg(dcache_n_161),
        .doUncachedResp_reg_0(dcache_n_580),
        .frontend_io_ptw_ptbr_mode(frontend_io_ptw_ptbr_mode),
        .frontend_io_ptw_req_ready(frontend_io_ptw_req_ready),
        .frontend_io_ptw_status_prv(frontend_io_ptw_status_prv[1]),
        .host_clk(host_clk),
        .invalid_paddr(invalid_paddr),
        .io_enq_bits_address(tlMasterXbar_auto_out_c_bits_address[11:6]),
        .lastGrant(\arb/lastGrant ),
        .lastGrant_reg(frontend_n_44),
        .pte_v(pte_v),
        .r_pte_d(r_pte_d),
        .\r_pte_ppn_reg[19]_0 (ptw_n_52),
        .\r_pte_ppn_reg[4]_0 (core_n_1800),
        .\r_pte_ppn_reg[4]_1 (core_n_1802),
        .\r_pte_ppn_reg[4]_2 (core_n_1804),
        .\r_pte_ppn_reg[4]_3 (core_n_1806),
        .\r_pte_ppn_reg[4]_4 (core_n_1809),
        .\r_pte_ppn_reg[4]_5 (core_n_1811),
        .\r_pte_ppn_reg[4]_6 (core_n_1813),
        .\r_pte_ppn_reg[4]_7 (core_n_1815),
        .r_pte_v_reg_0(dcache_n_582),
        .\r_refill_tag_reg[26] (arb_io_out_bits_addr),
        .\r_refill_waddr_reg[0] (ptw_n_73),
        .\reg_entries_0_reg[0] (ptw_n_134),
        .\reg_entries_0_reg[0]_0 ({ptw_n_135,ptw_n_136}),
        .\reg_entries_0_reg[0]_1 (ptw_n_160),
        .\reg_entries_0_reg[0]_10 (ptw_n_177),
        .\reg_entries_0_reg[0]_11 (ptw_n_178),
        .\reg_entries_0_reg[0]_12 (ptw_n_182),
        .\reg_entries_0_reg[0]_13 (ptw_n_183),
        .\reg_entries_0_reg[0]_14 (ptw_n_193),
        .\reg_entries_0_reg[0]_15 (\tlb/_T_210 ),
        .\reg_entries_0_reg[0]_16 (ptw_n_195),
        .\reg_entries_0_reg[0]_17 (ptw_n_196),
        .\reg_entries_0_reg[0]_18 (ptw_n_197),
        .\reg_entries_0_reg[0]_19 (\tlb/_T_194 ),
        .\reg_entries_0_reg[0]_2 (ptw_n_163),
        .\reg_entries_0_reg[0]_3 ({ptw_n_164,ptw_n_165}),
        .\reg_entries_0_reg[0]_4 (ptw_n_167),
        .\reg_entries_0_reg[0]_5 (ptw_n_168),
        .\reg_entries_0_reg[0]_6 (ptw_n_170),
        .\reg_entries_0_reg[0]_7 (ptw_n_172),
        .\reg_entries_0_reg[0]_8 (ptw_n_174),
        .\reg_entries_0_reg[0]_9 (ptw_n_176),
        .\reg_entries_0_reg[12] ({dcache_io_ptw_resp_bits_pte_u,dcache_io_ptw_resp_bits_pte_g,dcache_io_ptw_resp_bits_ae,\tlb/_T_943_4 }),
        .\reg_entries_0_reg[1] ({ptw_n_186,ptw_n_187}),
        .\reg_entries_0_reg[1]_0 ({ptw_n_188,ptw_n_189}),
        .\reg_entries_0_reg[1]_1 (\tlb/_T_728 ),
        .\reg_entries_0_reg[2] (\tlb/_T_382_3 ),
        .\reg_entries_0_reg[2]_0 (ptw_n_161),
        .\reg_entries_0_reg[2]_1 (ptw_n_166),
        .\reg_entries_0_reg[2]_2 (ptw_n_185),
        .\reg_entries_0_reg[2]_3 (\tlb/_T_482 ),
        .\reg_entries_0_reg[4] (ptw_n_15),
        .\reg_entries_0_reg[4]_0 (ptw_n_138),
        .\reg_entries_0_reg[4]_1 (ptw_n_148),
        .\reg_entries_0_reg[4]_2 (ptw_n_152),
        .\reg_entries_0_reg[4]_3 (ptw_n_154),
        .\reg_entries_0_reg[4]_4 (ptw_n_155),
        .\reg_entries_0_reg[4]_5 (ptw_n_156),
        .\reg_entries_0_reg[4]_6 (ptw_n_157),
        .\reg_entries_0_reg[4]_7 (ptw_n_159),
        .\reg_entries_0_reg[4]_8 (ptw_n_171),
        .\reg_entries_0_reg[4]_9 (ptw_n_180),
        .\reg_entries_0_reg[5] (ptw_n_53),
        .\reg_entries_0_reg[5]_0 (\tlb/_T_384 ),
        .\reg_entries_0_reg[6] (ptw_n_13),
        .\reg_entries_0_reg[6]_0 (ptw_n_14),
        .\reg_entries_0_reg[6]_1 (ptw_n_137),
        .\reg_entries_0_reg[6]_10 (ptw_n_147),
        .\reg_entries_0_reg[6]_11 (ptw_n_149),
        .\reg_entries_0_reg[6]_12 ({ptw_n_150,ptw_n_151}),
        .\reg_entries_0_reg[6]_13 (ptw_n_153),
        .\reg_entries_0_reg[6]_14 (ptw_n_158),
        .\reg_entries_0_reg[6]_15 (ptw_n_162),
        .\reg_entries_0_reg[6]_16 (ptw_n_169),
        .\reg_entries_0_reg[6]_17 (ptw_n_173),
        .\reg_entries_0_reg[6]_18 (ptw_n_175),
        .\reg_entries_0_reg[6]_19 (ptw_n_179),
        .\reg_entries_0_reg[6]_2 (ptw_n_139),
        .\reg_entries_0_reg[6]_20 (ptw_n_181),
        .\reg_entries_0_reg[6]_21 (ptw_n_184),
        .\reg_entries_0_reg[6]_22 (ptw_n_191),
        .\reg_entries_0_reg[6]_23 (ptw_n_192),
        .\reg_entries_0_reg[6]_24 (\tlb/_T_392 ),
        .\reg_entries_0_reg[6]_3 (ptw_n_140),
        .\reg_entries_0_reg[6]_4 (ptw_n_141),
        .\reg_entries_0_reg[6]_5 (ptw_n_142),
        .\reg_entries_0_reg[6]_6 (ptw_n_143),
        .\reg_entries_0_reg[6]_7 (ptw_n_144),
        .\reg_entries_0_reg[6]_8 (ptw_n_145),
        .\reg_entries_0_reg[6]_9 (ptw_n_146),
        .\reg_entries_0_reg[9] ({\tlb/_T_936 ,\tlb/_T_943 ,\tlb/_T_928 }),
        .\reg_entries_1_reg[0] (ptw_n_77),
        .\reg_entries_1_reg[0]_0 (ptw_n_85),
        .\reg_entries_1_reg[0]_1 (ptw_n_86),
        .\reg_entries_1_reg[0]_10 (ptw_n_95),
        .\reg_entries_1_reg[0]_11 (ptw_n_96),
        .\reg_entries_1_reg[0]_12 (ptw_n_97),
        .\reg_entries_1_reg[0]_13 (ptw_n_98),
        .\reg_entries_1_reg[0]_14 (ptw_n_99),
        .\reg_entries_1_reg[0]_15 (ptw_n_100),
        .\reg_entries_1_reg[0]_16 (ptw_n_101),
        .\reg_entries_1_reg[0]_17 (ptw_n_102),
        .\reg_entries_1_reg[0]_18 (ptw_n_104),
        .\reg_entries_1_reg[0]_19 (ptw_n_105),
        .\reg_entries_1_reg[0]_2 (ptw_n_87),
        .\reg_entries_1_reg[0]_20 (ptw_n_106),
        .\reg_entries_1_reg[0]_21 (ptw_n_107),
        .\reg_entries_1_reg[0]_22 (ptw_n_109),
        .\reg_entries_1_reg[0]_23 (ptw_n_110),
        .\reg_entries_1_reg[0]_24 (ptw_n_111),
        .\reg_entries_1_reg[0]_25 (ptw_n_112),
        .\reg_entries_1_reg[0]_26 (ptw_n_113),
        .\reg_entries_1_reg[0]_27 (ptw_n_114),
        .\reg_entries_1_reg[0]_28 (ptw_n_115),
        .\reg_entries_1_reg[0]_29 (ptw_n_116),
        .\reg_entries_1_reg[0]_3 (ptw_n_88),
        .\reg_entries_1_reg[0]_30 (ptw_n_117),
        .\reg_entries_1_reg[0]_31 (ptw_n_118),
        .\reg_entries_1_reg[0]_32 (ptw_n_119),
        .\reg_entries_1_reg[0]_33 (ptw_n_120),
        .\reg_entries_1_reg[0]_34 (ptw_n_121),
        .\reg_entries_1_reg[0]_35 (ptw_n_122),
        .\reg_entries_1_reg[0]_36 (_T_1488),
        .\reg_entries_1_reg[0]_37 (_T_1413),
        .\reg_entries_1_reg[0]_38 (_T_1338),
        .\reg_entries_1_reg[0]_39 (_T_1263),
        .\reg_entries_1_reg[0]_4 (ptw_n_89),
        .\reg_entries_1_reg[0]_40 (_T_1188),
        .\reg_entries_1_reg[0]_41 (_T_963),
        .\reg_entries_1_reg[0]_42 (_T_1113),
        .\reg_entries_1_reg[0]_43 (_T_1038),
        .\reg_entries_1_reg[0]_5 (ptw_n_90),
        .\reg_entries_1_reg[0]_6 (ptw_n_91),
        .\reg_entries_1_reg[0]_7 (ptw_n_92),
        .\reg_entries_1_reg[0]_8 (ptw_n_93),
        .\reg_entries_1_reg[0]_9 (ptw_n_94),
        .\reg_entries_4_reg[61] ({\tlb/p_0_in_1 [19],\tlb/p_0_in_1 [16],\tlb/p_0_in_1 [13]}),
        .\reg_entries_4_reg[61]_0 (\tlb/p_0_in ),
        .\reg_entries_4_reg[61]_1 (dcache_n_642),
        .\reg_entries_4_reg[61]_2 (dcache_n_643),
        .\reg_pmp_0_addr_reg[10] (core_n_518),
        .\reg_pmp_0_addr_reg[22] (core_n_1812),
        .\reg_pmp_0_addr_reg[28] (core_n_646),
        .\reg_pmp_0_addr_reg[28]_0 (core_n_1830),
        .\reg_pmp_0_addr_reg[28]_1 (core_n_1829),
        .\reg_pmp_0_addr_reg[29] ({frontend_io_ptw_pmp_0_addr[29:9],frontend_io_ptw_pmp_0_addr[0]}),
        .\reg_pmp_0_addr_reg[29]_0 (dcache_n_622),
        .\reg_pmp_1_addr_reg[22] (core_n_1816),
        .\reg_pmp_1_addr_reg[22]_0 (core_n_2006),
        .\reg_pmp_1_addr_reg[26] ({frontend_io_ptw_pmp_1_mask[29],frontend_io_ptw_pmp_1_mask[20],frontend_io_ptw_pmp_1_mask[11]}),
        .\reg_pmp_1_addr_reg[28] (core_n_645),
        .\reg_pmp_1_addr_reg[28]_0 (core_n_1832),
        .\reg_pmp_1_addr_reg[28]_1 (core_n_1831),
        .\reg_pmp_1_addr_reg[28]_2 (core_n_2004),
        .\reg_pmp_1_addr_reg[29] ({frontend_io_ptw_pmp_1_addr[29],frontend_io_ptw_pmp_1_addr[27:9],frontend_io_ptw_pmp_1_addr[0]}),
        .\reg_pmp_2_addr_reg[10] (core_n_519),
        .\reg_pmp_2_addr_reg[22] (core_n_1814),
        .\reg_pmp_2_addr_reg[26] ({frontend_io_ptw_pmp_2_mask[29],frontend_io_ptw_pmp_2_mask[20],frontend_io_ptw_pmp_2_mask[11]}),
        .\reg_pmp_2_addr_reg[28] (core_n_641),
        .\reg_pmp_2_addr_reg[28]_0 (core_n_1821),
        .\reg_pmp_2_addr_reg[28]_1 (core_n_1822),
        .\reg_pmp_2_addr_reg[29] ({frontend_io_ptw_pmp_2_addr[29:9],frontend_io_ptw_pmp_2_addr[0]}),
        .\reg_pmp_2_addr_reg[29]_0 (dcache_n_618),
        .\reg_pmp_3_addr_reg[22] (core_n_1810),
        .\reg_pmp_3_addr_reg[24] (core_n_459),
        .\reg_pmp_3_addr_reg[28] (core_n_640),
        .\reg_pmp_3_addr_reg[28]_0 (core_n_1819),
        .\reg_pmp_3_addr_reg[28]_1 (core_n_1820),
        .\reg_pmp_3_addr_reg[29] ({frontend_io_ptw_pmp_3_addr[29],frontend_io_ptw_pmp_3_addr[27:10]}),
        .\reg_pmp_3_cfg_a_reg[1] (core_n_1808),
        .\reg_pmp_4_addr_reg[10] (core_n_520),
        .\reg_pmp_4_addr_reg[22] (core_n_1807),
        .\reg_pmp_4_addr_reg[26] ({frontend_io_ptw_pmp_4_mask[29],frontend_io_ptw_pmp_4_mask[20],frontend_io_ptw_pmp_4_mask[11]}),
        .\reg_pmp_4_addr_reg[28] (core_n_639),
        .\reg_pmp_4_addr_reg[28]_0 (core_n_1817),
        .\reg_pmp_4_addr_reg[28]_1 (core_n_1818),
        .\reg_pmp_4_addr_reg[29] ({frontend_io_ptw_pmp_4_addr[29:9],frontend_io_ptw_pmp_4_addr[0]}),
        .\reg_pmp_4_addr_reg[29]_0 (dcache_n_620),
        .\reg_pmp_4_cfg_a_reg[1] (frontend_io_ptw_pmp_4_cfg_a),
        .\reg_pmp_5_addr_reg[22] (core_n_1805),
        .\reg_pmp_5_addr_reg[26] ({frontend_io_ptw_pmp_5_mask[29],frontend_io_ptw_pmp_5_mask[20],frontend_io_ptw_pmp_5_mask[11]}),
        .\reg_pmp_5_addr_reg[28] (core_n_642),
        .\reg_pmp_5_addr_reg[28]_0 (core_n_1823),
        .\reg_pmp_5_addr_reg[28]_1 (core_n_1824),
        .\reg_pmp_5_addr_reg[28]_2 (core_n_2005),
        .\reg_pmp_5_addr_reg[29] ({frontend_io_ptw_pmp_5_addr[29:9],frontend_io_ptw_pmp_5_addr[0]}),
        .\reg_pmp_5_cfg_a_reg[1] (frontend_io_ptw_pmp_5_cfg_a),
        .\reg_pmp_6_addr_reg[22] (core_n_1803),
        .\reg_pmp_6_addr_reg[26] ({frontend_io_ptw_pmp_6_mask[29],frontend_io_ptw_pmp_6_mask[20],frontend_io_ptw_pmp_6_mask[11]}),
        .\reg_pmp_6_addr_reg[28] (core_n_643),
        .\reg_pmp_6_addr_reg[28]_0 (core_n_1825),
        .\reg_pmp_6_addr_reg[28]_1 (core_n_1826),
        .\reg_pmp_6_addr_reg[28]_2 (core_n_2003),
        .\reg_pmp_6_addr_reg[29] ({frontend_io_ptw_pmp_6_addr[29:9],frontend_io_ptw_pmp_6_addr[0]}),
        .\reg_pmp_7_addr_reg[22] (core_n_1801),
        .\reg_pmp_7_addr_reg[24] (core_n_1927),
        .\reg_pmp_7_addr_reg[26] ({frontend_io_ptw_pmp_7_mask[29],frontend_io_ptw_pmp_7_mask[20],frontend_io_ptw_pmp_7_mask[11]}),
        .\reg_pmp_7_addr_reg[28] (core_n_644),
        .\reg_pmp_7_addr_reg[28]_0 (core_n_1827),
        .\reg_pmp_7_addr_reg[28]_1 (core_n_1828),
        .\reg_pmp_7_addr_reg[29] ({frontend_io_ptw_pmp_7_addr[29],frontend_io_ptw_pmp_7_addr[27:10]}),
        .\reg_sptbr_ppn_reg[19] (ptw_io_dpath_ptbr_ppn),
        .resp_valid_0_reg_0(dcache_n_635),
        .resp_valid_0_reg_1({dcache_n_636,dcache_n_637}),
        .resp_valid_0_reg_2(dcache_n_639),
        .resp_valid_0_reg_3(dcache_n_640),
        .resp_valid_0_reg_4(dcache_n_641),
        .resp_valid_0_reg_5({dcache_n_610,dcache_n_611}),
        .s0_clk_en(s0_clk_en),
        .\s1_pc_reg[28] (frontend_n_125),
        .\s1_pc_reg[31] ({s1_pc[31],s1_pc[28],s1_pc[25]}),
        .\s1_req_addr_reg[11] (core_n_1842),
        .\s1_req_addr_reg[11]_0 (core_n_1843),
        .\s1_req_addr_reg[32] ({dcache_n_139,dcache_n_140,dcache_n_141,dcache_n_142,dcache_n_143,dcache_n_144,dcache_n_145,dcache_n_146,dcache_n_147,dcache_n_148,dcache_n_149,dcache_n_150,dcache_n_151,dcache_n_152,dcache_n_153,dcache_n_154,dcache_n_155,dcache_n_156,dcache_n_157,dcache_n_158,dcache_n_159,_T_628}),
        .\s1_req_addr_reg[3] (dcache_n_631),
        .\s1_req_addr_reg[5] (dcache_n_625),
        .\s1_req_addr_reg[5]_0 (dcache_n_627),
        .\s1_req_addr_reg[7] (dcache_n_629),
        .\s1_req_addr_reg[7]_0 (dcache_n_628),
        .\s1_req_addr_reg[7]_1 (dcache_n_626),
        .\s1_req_addr_reg[7]_2 (dcache_n_632),
        .\s1_req_addr_reg[9] (dcache_n_630),
        .\s1_req_cmd_reg[4] (ptw_n_1),
        .\s1_req_cmd_reg[4]_0 (ptw_n_2),
        .\s1_req_cmd_reg[4]_1 (ptw_n_55),
        .s1_req_phys_reg(core_n_423),
        .s1_req_phys_reg_0(dcache_n_89),
        .s1_req_phys_reg_1(dcache_n_638),
        .s1_req_phys_reg_2(dcache_n_612),
        .s1_valid(s1_valid),
        .\s2_data_reg[10] (dcache_n_368),
        .\s2_data_reg[11] (dcache_n_370),
        .\s2_data_reg[12] (dcache_n_371),
        .\s2_data_reg[13] (dcache_n_372),
        .\s2_data_reg[14] (dcache_n_373),
        .\s2_data_reg[15] (dcache_n_374),
        .\s2_data_reg[16] (dcache_n_375),
        .\s2_data_reg[17] (dcache_n_376),
        .\s2_data_reg[18] (dcache_n_377),
        .\s2_data_reg[19] (dcache_n_378),
        .\s2_data_reg[20] (dcache_n_379),
        .\s2_data_reg[21] (dcache_n_380),
        .\s2_data_reg[22] (dcache_n_381),
        .\s2_data_reg[23] (dcache_n_382),
        .\s2_data_reg[24] (dcache_n_383),
        .\s2_data_reg[25] (dcache_n_384),
        .\s2_data_reg[26] (dcache_n_385),
        .\s2_data_reg[27] (dcache_n_386),
        .\s2_data_reg[28] (dcache_n_387),
        .\s2_data_reg[29] (dcache_n_388),
        .\s2_req_addr_reg[0] (dcache_n_443),
        .\s2_req_addr_reg[0]_0 (dcache_n_442),
        .\s2_req_addr_reg[0]_1 (dcache_n_441),
        .\s2_req_addr_reg[0]_2 (dcache_n_440),
        .\s2_req_addr_reg[0]_3 (dcache_n_439),
        .\s2_req_addr_reg[0]_4 (dcache_n_438),
        .\s2_req_cmd_reg[1] (dcache_n_583),
        .\s2_req_typ_reg[0] (dcache_n_567),
        .\s2_req_typ_reg[0]_0 (dcache_n_569),
        .\s2_req_typ_reg[0]_1 (dcache_n_570),
        .\s2_req_typ_reg[0]_2 (dcache_n_571),
        .\s2_req_typ_reg[0]_3 (dcache_n_572),
        .\s2_req_typ_reg[0]_4 (dcache_n_573),
        .\s2_req_typ_reg[0]_5 (dcache_n_574),
        .\s2_req_typ_reg[0]_6 (dcache_n_575),
        .\s2_req_typ_reg[0]_7 (dcache_n_367),
        .s2_valid_reg(s2_valid_reg),
        .state(\tlb/state_2 ),
        .state_0(\tlb/state ),
        .\state_reg[0]_0 (ptw_n_16),
        .\state_reg[0]_1 (ptw_n_131),
        .\state_reg[0]_2 (dcache_n_576),
        .\state_reg[1]_0 (ptw_n_37),
        .\state_reg[1]_1 (ptw_n_72),
        .target_reset(target_reset),
        .traverse(traverse),
        .\valid_reg[3] (ptw_n_132));
  LUT1 #(
    .INIT(2'h1)) 
    \remainder[103]_i_13 
       (.I0(core_n_357),
        .O(\remainder[103]_i_13_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \remainder[103]_i_14 
       (.I0(core_n_357),
        .O(\remainder[103]_i_14_n_0 ));
  CARRY4 \s1_pc_reg[39]_i_10 
       (.CI(\s1_pc_reg[39]_i_12_n_0 ),
        .CO(_T_2181),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,core_n_651}));
  CARRY4 \s1_pc_reg[39]_i_11 
       (.CI(\s1_pc_reg[39]_i_14_n_0 ),
        .CO(_T_2179),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,core_n_1705}));
  CARRY4 \s1_pc_reg[39]_i_12 
       (.CI(\s1_pc_reg[39]_i_16_n_0 ),
        .CO({\s1_pc_reg[39]_i_12_n_0 ,\s1_pc_reg[39]_i_12_n_1 ,\s1_pc_reg[39]_i_12_n_2 ,\s1_pc_reg[39]_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1434,core_n_1435,core_n_1436,core_n_1437}));
  CARRY4 \s1_pc_reg[39]_i_14 
       (.CI(\s1_pc_reg[39]_i_21_n_0 ),
        .CO({\s1_pc_reg[39]_i_14_n_0 ,\s1_pc_reg[39]_i_14_n_1 ,\s1_pc_reg[39]_i_14_n_2 ,\s1_pc_reg[39]_i_14_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1442,core_n_1443,core_n_1444,core_n_1445}));
  CARRY4 \s1_pc_reg[39]_i_16 
       (.CI(\<const0> ),
        .CO({\s1_pc_reg[39]_i_16_n_0 ,\s1_pc_reg[39]_i_16_n_1 ,\s1_pc_reg[39]_i_16_n_2 ,\s1_pc_reg[39]_i_16_n_3 }),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1430,core_n_1431,core_n_1432,core_n_1433}));
  CARRY4 \s1_pc_reg[39]_i_21 
       (.CI(\<const0> ),
        .CO({\s1_pc_reg[39]_i_21_n_0 ,\s1_pc_reg[39]_i_21_n_1 ,\s1_pc_reg[39]_i_21_n_2 ,\s1_pc_reg[39]_i_21_n_3 }),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1438,core_n_1439,core_n_1440,core_n_1441}));
  CARRY4 \s1_req_addr_reg[39]_i_13 
       (.CI(\<const0> ),
        .CO({\s1_req_addr_reg[39]_i_13_n_0 ,\s1_req_addr_reg[39]_i_13_n_1 ,\s1_req_addr_reg[39]_i_13_n_2 ,\s1_req_addr_reg[39]_i_13_n_3 }),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1612,core_n_1613,core_n_1614,core_n_1615}));
  CARRY4 \s1_req_addr_reg[39]_i_2 
       (.CI(\s1_req_addr_reg[39]_i_4_n_0 ),
        .CO(_T_2774),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,_T_2770[24]}));
  CARRY4 \s1_req_addr_reg[39]_i_3 
       (.CI(\s1_req_addr_reg[39]_i_6_n_0 ),
        .CO(_T_2772),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,\<const0> ,core_n_1787}));
  CARRY4 \s1_req_addr_reg[39]_i_4 
       (.CI(\s1_req_addr_reg[39]_i_8_n_0 ),
        .CO({\s1_req_addr_reg[39]_i_4_n_0 ,\s1_req_addr_reg[39]_i_4_n_1 ,\s1_req_addr_reg[39]_i_4_n_2 ,\s1_req_addr_reg[39]_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1688,core_n_1689,core_n_1690,core_n_1691}));
  CARRY4 \s1_req_addr_reg[39]_i_6 
       (.CI(\s1_req_addr_reg[39]_i_13_n_0 ),
        .CO({\s1_req_addr_reg[39]_i_6_n_0 ,\s1_req_addr_reg[39]_i_6_n_1 ,\s1_req_addr_reg[39]_i_6_n_2 ,\s1_req_addr_reg[39]_i_6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1692,core_n_1693,core_n_1694,core_n_1695}));
  CARRY4 \s1_req_addr_reg[39]_i_8 
       (.CI(\<const0> ),
        .CO({\s1_req_addr_reg[39]_i_8_n_0 ,\s1_req_addr_reg[39]_i_8_n_1 ,\s1_req_addr_reg[39]_i_8_n_2 ,\s1_req_addr_reg[39]_i_8_n_3 }),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1608,core_n_1609,core_n_1610,core_n_1611}));
  TLBuffer_19 sync_xing
       (.ADDRARDADDR({sync_xing_n_54,sync_xing_n_55,sync_xing_n_56,sync_xing_n_57,sync_xing_n_58,sync_xing_n_59}),
        .ADDRBWRADDR(ADDRBWRADDR[0]),
        .CO(\_T_5874_reg[0] ),
        .DIA(tlMasterXbar_auto_out_c_bits_size),
        .DIB(tlMasterXbar_auto_out_a_bits_opcode),
        .DOA(sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_opcode[1:0]),
        .DOB(sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_opcode[2]),
        .DOBDO({dcache_n_0,dcache_n_1,dcache_n_2,dcache_n_3,dcache_n_4,dcache_n_5,dcache_n_6,dcache_n_7}),
        .E(sync_xing_n_41),
        .SR(sync_xing_n_365),
        .WEBWE(sync_xing_n_40),
        .\_T_1052_reg[0] (tlMasterXbar_n_7),
        .\_T_1052_reg[7] (sync_xing_n_49),
        ._T_1053_reg(_T_1053_reg),
        .\_T_1055_reg[25] (io_enq_bits_address),
        .\_T_1057_reg[0] (\_T_1057_reg[0] ),
        .\_T_1057_reg[0]_0 (\_T_1057_reg[0]_0 ),
        .\_T_1057_reg[1] (\_T_1057_reg[1] ),
        .\_T_1057_reg[1]_0 (\_T_1057_reg[1]_0 ),
        .\_T_1057_reg[1]_1 (\_T_1057_reg[1]_1 ),
        .\_T_1066_reg[0] (sync_xing_n_366),
        .\_T_1066_reg[0]_0 (tlMasterXbar_n_4),
        .\_T_1066_reg[1] (tlMasterXbar_n_5),
        ._T_1161_1(_T_1161_1),
        ._T_1172_1(_T_1172_1),
        ._T_1208({_T_1208[114:110],_T_1208[106],_T_1208[104],_T_1208[77:72],_T_1208[63:0]}),
        .\_T_1250_reg[2] (\_T_1250_reg[2] ),
        ._T_1402(_T_1402),
        ._T_1567_reg(dcache_n_432),
        ._T_1670_reg(_T_1670_reg),
        .\_T_191_reg[0] (\icache/_T_191_reg__0 ),
        .\_T_191_reg[1] (sync_xing_n_43),
        .\_T_191_reg[2] (sync_xing_n_42),
        .\_T_191_reg[3] (sync_xing_n_44),
        .\_T_191_reg[3]_0 (frontend_n_244),
        .\_T_191_reg[3]_1 (frontend_n_240),
        .\_T_191_reg[5] (sync_xing_n_46),
        .\_T_191_reg[5]_0 (frontend_n_243),
        .\_T_191_reg[7] (sync_xing_n_47),
        .\_T_191_reg[7]_0 (frontend_n_241),
        .\_T_191_reg[8] (tlMasterXbar_auto_in_0_d_bits_size),
        .\_T_191_reg[8]_0 ({\icache/p_0_in__0 [8],\icache/p_0_in__0 [6],\icache/p_0_in__0 [4],\icache/p_0_in__0 [0]}),
        .\_T_191_reg[8]_1 (frontend_n_245),
        .\_T_250_0_bits_data_reg[61] (ram_data__T_63_data),
        .\_T_3585_reg[0] (p_0_in_5),
        .\_T_3585_reg[1] (sync_xing_n_356),
        .\_T_3585_reg[1]_0 (_T_3585_reg__0),
        .\_T_3585_reg[2] (dcache_n_415),
        .\_T_3585_reg[3] (sync_xing_n_354),
        .\_T_3585_reg[5] (sync_xing_n_357),
        .\_T_3585_reg[5]_0 (dcache_n_448),
        .\_T_3585_reg[6] (sync_xing_n_352),
        .\_T_3585_reg[6]_0 (dcache_n_453),
        .\_T_3585_reg[7] (sync_xing_n_358),
        .\_T_3585_reg[7]_0 (dcache_n_454),
        ._T_3628(_T_3628),
        .\_T_3859_reg[8] (sync_xing_n_22),
        .\_T_4992_reg[2] (\_T_4992_reg[2] ),
        .\_T_4992_reg[3] (\_T_4992_reg[3] ),
        .\_T_4992_reg[6] (\_T_4992_reg[6] ),
        .\_T_4992_reg[7] (\_T_4992_reg[7] ),
        .\_T_4992_reg[8] (\_T_4992_reg[8] ),
        .\_T_5010_reg[1] (\_T_5010_reg[1] ),
        ._T_5195_0_reg(_T_5195_0_reg),
        .\_T_5351_reg[0] (sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_size[3:2]),
        .\_T_5351_reg[0]_0 (\_T_5351_reg[0] ),
        .\_T_5351_reg[0]_1 (\_T_5351_reg[0]_0 ),
        .\_T_5351_reg[3] (\_T_5351_reg[3] ),
        .\_T_5369_reg[1] (\_T_5369_reg[1] ),
        .\_T_5369_reg[5] (\_T_5369_reg[5] ),
        ._T_5554_4_reg(_T_5554_4_reg),
        ._T_5577_0(_T_5577_0),
        .\_T_558_reg[2] (\_T_558_reg[2] ),
        .\_T_5856_reg[0] (\_T_5856_reg[0] ),
        .\_T_5856_reg[1] (\_T_5856_reg[1] ),
        .\_T_5856_reg[2] (\_T_5856_reg[2] ),
        .\_T_5856_reg[3] (\_T_5856_reg[3] ),
        .\_T_5856_reg[5] (\_T_5856_reg[5] ),
        .\_T_5874_reg[1] (\_T_5874_reg[1] ),
        .\_T_5874_reg[1]_0 (sbus_auto_coupler_from_tile_named_tile_fixer_in_a_valid),
        .\_T_5874_reg[1]_1 (\_T_5874_reg[1]_0 ),
        .\_T_5874_reg[2] (\_T_5874_reg[2] ),
        ._T_6059_0_reg(_T_6059_0_reg),
        .\_T_6215_reg[1] (\_T_6215_reg[1] ),
        .\_T_6215_reg[2] (\_T_6215_reg[2] ),
        .\_T_6215_reg[3] (\_T_6215_reg[3] ),
        .\_T_6233_reg[0] (\_T_6233_reg[0] ),
        .\_T_6233_reg[0]_0 (\_T_6233_reg[0]_0 ),
        .\_T_6233_reg[1] (\_T_6233_reg[1] ),
        .\_T_6233_reg[1]_0 (\_T_6233_reg[1]_0 ),
        .\_T_6233_reg[5] (\_T_6233_reg[5] ),
        .\_T_6233_reg[5]_0 (\_T_6233_reg[5]_0 ),
        .\_T_6233_reg[5]_1 (\_T_6233_reg[5]_1 ),
        ._T_6418_0_reg(_T_6418_0_reg),
        ._T_642_0(_T_642_0),
        ._T_642_1_reg(_T_642_1_reg),
        .\_T_6648_reg[2] (\_T_6648_reg[2] ),
        ._T_6804_0_reg(_T_6804_0_reg),
        .\_T_767_reg[0] (sbus_auto_coupler_to_mbus_nodelay_out_c_bits_size[2]),
        .\_T_767_reg[2] (\_T_767_reg[2] ),
        .\_T_767_reg[2]_0 (\_T_767_reg[2]_0 ),
        ._T_920_0(_T_920_0),
        ._T_920_0_reg(_T_920_0_reg),
        ._T_920_1(_T_920_1),
        ._T_920_1_reg(_T_920_1_reg),
        ._T_920_3_reg(_T_920_3_reg),
        ._T_940_0(_T_940_0),
        .\address_reg[30] (\address_reg[30] ),
        .\address_reg[31] (\address_reg[31] ),
        .\address_reg[31]_0 (\address_reg[31]_0 ),
        .\address_reg[31]_1 (\address_reg[31]_1 ),
        .\address_reg[31]_2 (\address_reg[31]_2 ),
        .\beatsLeft_reg[1] (\beatsLeft_reg[1] ),
        .bh_auto_out_a_ready(bh_auto_out_a_ready),
        .blockProbeAfterGrantCount(blockProbeAfterGrantCount),
        .blockUncachedGrant(blockUncachedGrant),
        .count_reg(count_reg),
        .count_reg_0(count_reg_0),
        .count_reg_1(count_reg_1),
        .count_reg_2(count_reg_2),
        .count_reg_3(count_reg_3),
        .count_reg_4(count_reg_4),
        .count_reg_5(count_reg_5),
        .count_reg_6(count_reg_6),
        .count_reg_7(count_reg_7),
        .count_reg_8(count_reg_8),
        .dataArb_io_in_1_valid(dataArb_io_in_1_valid),
        .data_arrays_0_0_reg(tlMasterXbar_auto_in_0_d_bits_opcode),
        .data_arrays_0_0_reg_0(sync_xing_n_45),
        .data_arrays_0_0_reg_1(sync_xing_n_48),
        .data_arrays_0_0_reg_10(sync_xing_n_355),
        .data_arrays_0_0_reg_2(sync_xing_n_210),
        .data_arrays_0_0_reg_3(sync_xing_n_212),
        .data_arrays_0_0_reg_4(sync_xing_n_213),
        .data_arrays_0_0_reg_5(sync_xing_n_214),
        .data_arrays_0_0_reg_6(sync_xing_n_215),
        .data_arrays_0_0_reg_7(sync_xing_n_216),
        .data_arrays_0_0_reg_8(sync_xing_n_217),
        .data_arrays_0_0_reg_9(sync_xing_n_218),
        .data_arrays_0_1_reg({dcache_n_17,dcache_n_18,dcache_n_19,dcache_n_20,dcache_n_21,dcache_n_22,dcache_n_23,dcache_n_24}),
        .data_arrays_0_2_reg({dcache_n_25,dcache_n_26,dcache_n_27,dcache_n_28,dcache_n_29,dcache_n_30,dcache_n_31,dcache_n_32}),
        .data_arrays_0_3_reg({dcache_n_33,dcache_n_34,dcache_n_35,dcache_n_36,dcache_n_37,dcache_n_38,dcache_n_39,dcache_n_40}),
        .data_arrays_0_4_reg({dcache_n_41,dcache_n_42,dcache_n_43,dcache_n_44,dcache_n_45,dcache_n_46,dcache_n_47,dcache_n_48}),
        .data_arrays_0_5_reg({dcache_n_49,dcache_n_50,dcache_n_51,dcache_n_52,dcache_n_53,dcache_n_54,dcache_n_55,dcache_n_56}),
        .data_arrays_0_6_reg({dcache_n_57,dcache_n_58,dcache_n_59,dcache_n_60,dcache_n_61,dcache_n_62,dcache_n_63,dcache_n_64}),
        .data_arrays_0_7_reg(sync_xing_n_34),
        .data_arrays_0_7_reg_0({dcache_n_65,dcache_n_66,dcache_n_67,dcache_n_68,dcache_n_69,dcache_n_70,dcache_n_71,dcache_n_72}),
        .data_arrays_1_0_reg(sync_xing_n_35),
        .dcacheArb_io_requestor_1_replay_next(dcacheArb_io_requestor_1_replay_next),
        .got_e_reg(DOA),
        .got_e_reg_0(got_e_reg),
        .got_e_reg_1(got_e_reg_0),
        .grantInProgress_reg(sync_xing_n_51),
        .grantInProgress_reg_0(dcache_n_416),
        .grantInProgress_reg_1(dcache_n_75),
        .host_clk(host_clk),
        .invalidated(\icache/invalidated ),
        .io_enq_bits_address(tlMasterXbar_auto_out_a_bits_address),
        .io_enq_bits_data(io_enq_bits_data),
        .io_enq_bits_mask(tlMasterXbar_auto_out_a_bits_mask),
        .io_enq_bits_param(io_enq_bits_param),
        .io_enq_bits_source(io_enq_bits_source),
        .io_mask(fq_io_mask),
        .load(\icache/load ),
        .maybe_full(\Queue/maybe_full ),
        .maybe_full_3(\Queue_3/maybe_full ),
        .maybe_full_reg(maybe_full_reg),
        .maybe_full_reg_0(maybe_full_reg_0),
        .maybe_full_reg_1(maybe_full_reg_1),
        .mem_reg_valid_reg(mem_reg_replay_reg),
        .p_12_in(\icache/p_12_in ),
        .p_1_in(\Queue/p_1_in ),
        .\param_reg[1] (sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_param[1:0]),
        .\param_reg[2] (sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_param[2]),
        .\probe_bits_address_reg[10] (ptw_n_69),
        .\probe_bits_address_reg[11] (ptw_n_70),
        .\probe_bits_address_reg[31] (tlMasterXbar_auto_out_c_bits_address),
        .\probe_bits_address_reg[3] (dcache_n_417),
        .\probe_bits_address_reg[4] (dcache_n_418),
        .\probe_bits_address_reg[6] (ptw_n_56),
        .\probe_bits_address_reg[7] (ptw_n_66),
        .\probe_bits_address_reg[8] (ptw_n_67),
        .\probe_bits_address_reg[9] (ptw_n_68),
        .\probe_bits_param_reg[1] (_T_258),
        .\probe_bits_param_reg[1]_0 (sync_xing_n_220),
        .\probe_bits_size_reg[3] (tlMasterXbar_auto_in_0_b_bits_size),
        .probe_bits_source_reg(tlMasterXbar_auto_out_c_bits_source),
        .pstore1_rmw_reg(dcache_n_136),
        .pstore2_valid_reg(dcache_n_212),
        .ram_address__T_63_data(ram_address__T_63_data),
        .ram_data__T_63_data(tlMasterXbar_auto_in_0_d_bits_data),
        .\ram_data_reg[63] (\ram_data_reg[63] ),
        .\ram_id_reg[0] (\ram_id_reg[0] ),
        .\ram_id_reg[3] (\ram_id_reg[3] ),
        .\ram_id_reg[4] (\ram_id_reg[4] ),
        .\ram_id_reg[5] (\ram_id_reg[5] ),
        .ram_mask__T_63_data(ram_mask__T_63_data),
        .\ram_opcode_reg[1] (\ram_opcode_reg[1] ),
        .ram_param__T_63_data(tlMasterXbar_auto_in_0_b_bits_param),
        .\ram_size_reg[1] (DIB),
        .ram_source__T_63_data(ram_source__T_63_data),
        .\ram_strb_reg[0] (\ram_strb_reg[0] ),
        .\ram_strb_reg[0]_0 (\ram_strb_reg[0]_0 ),
        .\ram_strb_reg[1] (\ram_strb_reg[1] ),
        .\ram_strb_reg[2] (\ram_strb_reg[2] ),
        .\ram_strb_reg[2]_0 (\ram_strb_reg[2]_0 ),
        .\ram_strb_reg[3] (\ram_strb_reg[3] ),
        .\ram_strb_reg[4] (\ram_strb_reg[4] ),
        .\ram_strb_reg[4]_0 (\ram_strb_reg[4]_0 ),
        .\ram_strb_reg[5] (\ram_strb_reg[5] ),
        .\ram_strb_reg[6] (\ram_strb_reg[6] ),
        .\ram_strb_reg[6]_0 (\ram_strb_reg[6]_0 ),
        .\ram_strb_reg[7] (\ram_strb_reg[7] ),
        .\ram_user_reg[6] (\ram_user_reg[6] ),
        .\ram_user_reg[8] (sbus_auto_coupler_to_mbus_nodelay_out_c_bits_size[1:0]),
        .refill_one_beat(\icache/refill_one_beat ),
        .refill_valid_reg(sync_xing_n_33),
        .release_ack_wait30_out(release_ack_wait30_out),
        .release_ack_wait_reg(sync_xing_n_207),
        .release_ack_wait_reg_0(dcache_n_90),
        .\release_state_reg[0] (dcache_n_433),
        .\release_state_reg[1] (tlMasterXbar_auto_out_c_bits_opcode),
        .\release_state_reg[1]_0 ({dcache_n_137,dcache_n_138}),
        .resp_send_reg(resp_send_reg),
        .s1_probe_reg(sync_xing_n_359),
        .s1_release_data_valid(s1_release_data_valid),
        .s1_release_data_valid_reg(sync_xing_n_32),
        .\s1_req_addr_reg[31] (tlMasterXbar_auto_in_0_b_bits_address),
        .\s1_req_addr_reg[39] (sync_xing_n_50),
        .s1_valid(s1_valid),
        .s1_valid_reg(dcache_n_346),
        .\s2_data_reg[63] (_T_766),
        .\s2_data_reg[63]_0 (tlMasterXbar_auto_out_c_bits_data),
        .\s2_pc_reg[11] ({D,frontend_n_239}),
        .s2_release_data_valid0(s2_release_data_valid0),
        .\s2_req_addr_reg[10] ({_T_3959[10],_T_3959[8]}),
        .\s2_req_addr_reg[11] ({dataArb_io_in_1_bits_addr[11],dataArb_io_in_1_bits_addr[9],dataArb_io_in_1_bits_addr[7:6]}),
        .\s2_req_cmd_reg[0] (dcache_n_435),
        .\s2_req_cmd_reg[0]_0 (dcache_n_436),
        .\s2_req_cmd_reg[4] (dcache_n_213),
        .\saved_address_reg[1] (\saved_address_reg[1] ),
        .\saved_address_reg[1]_0 (\saved_address_reg[1]_0 ),
        .\saved_address_reg[7] (\saved_address_reg[7] ),
        .\saved_address_reg[7]_0 (\saved_address_reg[7]_0 ),
        .\saved_address_reg[7]_1 (\saved_address_reg[7]_1 ),
        .\saved_address_reg[7]_2 (\saved_address_reg[7]_2 ),
        .\saved_address_reg[7]_3 (\saved_address_reg[7]_3 ),
        .\saved_address_reg[7]_4 (\saved_address_reg[7]_4 ),
        .\saved_opcode_reg[1] (DIA),
        .sbus_auto_coupler_from_port_named_blkdevcontroller_passthru_in_0_a_bits_address(sbus_auto_coupler_from_port_named_blkdevcontroller_passthru_in_0_a_bits_address),
        .sbus_auto_coupler_from_port_named_blkdevcontroller_passthru_in_1_a_bits_address(sbus_auto_coupler_from_port_named_blkdevcontroller_passthru_in_1_a_bits_address),
        .sbus_auto_coupler_from_port_named_serialadapter_passthru_in_a_bits_address(sbus_auto_coupler_from_port_named_serialadapter_passthru_in_a_bits_address),
        .sbus_auto_coupler_from_port_named_serialadapter_passthru_in_a_bits_opcode(sbus_auto_coupler_from_port_named_serialadapter_passthru_in_a_bits_opcode),
        .sbus_auto_coupler_from_tile_named_tile_fixer_in_a_ready(sbus_auto_coupler_from_tile_named_tile_fixer_in_a_ready),
        .sbus_auto_coupler_from_tile_named_tile_fixer_in_b_valid(sbus_auto_coupler_from_tile_named_tile_fixer_in_b_valid),
        .sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_error(sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_error),
        .sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_opcode(sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_opcode),
        .sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_sink(sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_sink),
        .sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_size(sbus_auto_coupler_from_tile_named_tile_fixer_in_d_bits_size),
        .sbus_auto_coupler_from_tile_named_tile_fixer_in_d_ready(sbus_auto_coupler_from_tile_named_tile_fixer_in_d_ready),
        .sbus_auto_coupler_to_mbus_nodelay_out_a_bits_opcode(sbus_auto_coupler_to_mbus_nodelay_out_a_bits_opcode),
        .sbus_auto_coupler_to_mbus_nodelay_out_d_ready(sbus_auto_coupler_to_mbus_nodelay_out_d_ready),
        .\sendaddr_reg[11] (\sendaddr_reg[11] ),
        .\size_reg[1] (sbus_auto_coupler_from_tile_named_tile_fixer_in_a_bits_size[1:0]),
        .\source_reg[0] (\source_reg[0] ),
        .\source_reg[1] (\source_reg[1] ),
        .\source_reg[4] (\source_reg[4] ),
        .\state_reg[0] (\state_reg[0] ),
        .\state_reg[0]_0 (\state_reg[0]_0 ),
        .\state_reg[0]_1 (\state_reg[0]_1 ),
        .\state_reg[0]_2 (\state_reg[0]_2 ),
        .\state_reg[0]_3 (\state_reg[0]_3 ),
        .system_bus_xbar_auto_out_3_a_bits_param(system_bus_xbar_auto_out_3_a_bits_param),
        .tag_array_0_reg(sync_xing_n_208),
        .tag_array_0_reg_0(sync_xing_n_209),
        .tag_array_0_reg_1(dcache_n_423),
        .tag_array_0_reg_i_10__0(tag_array_0_reg_i_10__0),
        .tag_array_0_reg_i_11__0(tag_array_0_reg_i_11__0),
        .tag_array_0_reg_i_12__0(tag_array_0_reg_i_12__0),
        .tag_array_0_reg_i_13__0(tag_array_0_reg_i_13__0),
        .tag_array_0_reg_i_13__0_0(tag_array_0_reg_i_13__0_0),
        .tag_array_0_reg_i_8__0(tag_array_0_reg_i_8__0),
        .tag_array_0_reg_i_9__0(tag_array_0_reg_i_9__0),
        .target_reset(target_reset),
        .tlMasterXbar_auto_in_0_d_bits_error(tlMasterXbar_auto_in_0_d_bits_error),
        .tlMasterXbar_auto_out_a_bits_size(tlMasterXbar_auto_out_a_bits_size),
        .tlMasterXbar_auto_out_b_bits_source(tlMasterXbar_auto_out_b_bits_source),
        .uncachedInFlight_0_reg(sync_xing_n_350),
        .uncachedInFlight_0_reg_0(dcache_n_431),
        .value(\Queue/value ),
        .value_1(\Queue/value_1 ),
        .value_1_0(\Queue_3/value_1 ),
        .value_1_reg(value_1_reg),
        .\value_1_reg[0] (\value_1_reg[0] ),
        .\value_1_reg[1] (\value_1_reg[1] ),
        .value_2(\Queue_3/value ),
        .value_reg(tlMasterXbar_n_2),
        .value_reg_0(value_reg),
        .value_reg_1(value_reg_0),
        .\vb_array_reg[0] (sync_xing_n_39));
  TLXbar_5 tlMasterXbar
       (.DIB(tlMasterXbar_auto_out_a_bits_opcode),
        .Q(tlMasterXbar_auto_in_1_a_bits_address),
        .SR(sync_xing_n_365),
        .\_T_1052_reg[7]_0 (tlMasterXbar_n_5),
        .\_T_1066_reg[1]_0 (tlMasterXbar_n_7),
        ._T_1161_0_reg_0(tlMasterXbar_n_10),
        ._T_1161_1(_T_1161_1),
        ._T_1172_1(_T_1172_1),
        ._T_165_reg(frontend_n_49),
        .host_clk(host_clk),
        .io_enq_bits_address(tlMasterXbar_auto_out_a_bits_address),
        .io_enq_bits_mask(tlMasterXbar_auto_out_a_bits_mask[7:6]),
        .maybe_full(\Queue/maybe_full ),
        .maybe_full_reg(sync_xing_n_366),
        .p_1_in(\Queue/p_1_in ),
        .refill_valid_reg(tlMasterXbar_n_4),
        .release_ack_wait_reg(dcache_n_210),
        .release_ack_wait_reg_0(dcache_n_209),
        .\s2_req_addr_reg[31] ({_GEN_283_0,_T_3959}),
        .\s2_req_cmd_reg[4] (dcache_n_213),
        .s2_uncached(s2_uncached),
        .s2_uncached_reg(dcache_n_343),
        .s2_uncached_reg_0(dcache_n_455),
        .s2_uncached_reg_1(dcache_n_456),
        .s2_uncached_reg_2(dcache_n_342),
        .target_reset(target_reset),
        .tlMasterXbar_auto_in_0_a_bits_size(tlMasterXbar_auto_in_0_a_bits_size),
        .tlMasterXbar_auto_out_a_bits_size(tlMasterXbar_auto_out_a_bits_size[2]),
        .\uncachedReqs_0_addr_reg[2] (tlMasterXbar_n_6),
        .value(\Queue/value ),
        .value_1(\Queue/value_1 ),
        .value_reg(tlMasterXbar_n_2),
        .value_reg_0(sync_xing_n_49));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[11]_i_2 
       (.I0(core_n_1546),
        .I1(mem_reg_pc[11]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[24]),
        .O(\trig_pc[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[11]_i_3 
       (.I0(core_n_1547),
        .I1(mem_reg_pc[10]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[20]),
        .O(\trig_pc[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[11]_i_4 
       (.I0(core_n_1548),
        .I1(mem_reg_pc[9]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[19]),
        .O(\trig_pc[11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[11]_i_5 
       (.I0(core_n_1549),
        .I1(mem_reg_pc[8]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[18]),
        .O(\trig_pc[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[15]_i_2 
       (.I0(core_n_1542),
        .I1(mem_reg_pc[15]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[28]),
        .O(\trig_pc[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[15]_i_3 
       (.I0(core_n_1543),
        .I1(mem_reg_pc[14]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[27]),
        .O(\trig_pc[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[15]_i_4 
       (.I0(core_n_1544),
        .I1(mem_reg_pc[13]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[26]),
        .O(\trig_pc[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[15]_i_5 
       (.I0(core_n_1545),
        .I1(mem_reg_pc[12]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[25]),
        .O(\trig_pc[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[19]_i_2 
       (.I0(core_n_1538),
        .I1(mem_reg_pc[19]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[35]),
        .O(\trig_pc[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[19]_i_3 
       (.I0(core_n_1539),
        .I1(mem_reg_pc[18]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[34]),
        .O(\trig_pc[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[19]_i_4 
       (.I0(core_n_1540),
        .I1(mem_reg_pc[17]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[33]),
        .O(\trig_pc[19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[19]_i_5 
       (.I0(core_n_1541),
        .I1(mem_reg_pc[16]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[32]),
        .O(\trig_pc[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[23]_i_2 
       (.I0(core_n_1534),
        .I1(mem_reg_pc[23]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[42]),
        .O(\trig_pc[23]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[23]_i_3 
       (.I0(core_n_1535),
        .I1(mem_reg_pc[22]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[41]),
        .O(\trig_pc[23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[23]_i_4 
       (.I0(core_n_1536),
        .I1(mem_reg_pc[21]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[40]),
        .O(\trig_pc[23]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[23]_i_5 
       (.I0(core_n_1537),
        .I1(mem_reg_pc[20]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[36]),
        .O(\trig_pc[23]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[27]_i_2 
       (.I0(core_n_1530),
        .I1(mem_reg_pc[27]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[49]),
        .O(\trig_pc[27]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[27]_i_3 
       (.I0(core_n_1531),
        .I1(mem_reg_pc[26]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[48]),
        .O(\trig_pc[27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[27]_i_4 
       (.I0(core_n_1532),
        .I1(mem_reg_pc[25]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[44]),
        .O(\trig_pc[27]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[27]_i_5 
       (.I0(core_n_1533),
        .I1(mem_reg_pc[24]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[43]),
        .O(\trig_pc[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[31]_i_2 
       (.I0(core_n_1526),
        .I1(mem_reg_pc[31]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[56]),
        .O(\trig_pc[31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[31]_i_3 
       (.I0(core_n_1527),
        .I1(mem_reg_pc[30]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[52]),
        .O(\trig_pc[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[31]_i_4 
       (.I0(core_n_1528),
        .I1(mem_reg_pc[29]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[51]),
        .O(\trig_pc[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[31]_i_5 
       (.I0(core_n_1529),
        .I1(mem_reg_pc[28]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[50]),
        .O(\trig_pc[31]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[35]_i_2 
       (.I0(core_n_1522),
        .I1(mem_reg_pc[35]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[60]),
        .O(\trig_pc[35]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[35]_i_3 
       (.I0(core_n_1523),
        .I1(mem_reg_pc[34]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[59]),
        .O(\trig_pc[35]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[35]_i_4 
       (.I0(core_n_1524),
        .I1(mem_reg_pc[33]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[58]),
        .O(\trig_pc[35]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[35]_i_5 
       (.I0(core_n_1525),
        .I1(mem_reg_pc[32]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[57]),
        .O(\trig_pc[35]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[39]_i_2 
       (.I0(core_n_1518),
        .I1(mem_reg_pc[39]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[52]),
        .O(\trig_pc[39]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[39]_i_3 
       (.I0(core_n_1519),
        .I1(mem_reg_pc[38]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[52]),
        .O(\trig_pc[39]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[39]_i_4 
       (.I0(core_n_1520),
        .I1(mem_reg_pc[37]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[52]),
        .O(\trig_pc[39]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[39]_i_5 
       (.I0(core_n_1521),
        .I1(mem_reg_pc[36]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[52]),
        .O(\trig_pc[39]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[3]_i_2 
       (.I0(core_n_1554),
        .I1(mem_reg_pc[3]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[10]),
        .O(\trig_pc[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[3]_i_3 
       (.I0(core_n_1555),
        .I1(mem_reg_pc[2]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[9]),
        .O(\trig_pc[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[3]_i_4 
       (.I0(core_n_1556),
        .I1(mem_reg_pc[1]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[8]),
        .O(\trig_pc[3]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[43]_i_2 
       (.I0(core_n_1514),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[43]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[43]_i_3 
       (.I0(core_n_1515),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[43]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[43]_i_4 
       (.I0(core_n_1516),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[43]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[43]_i_5 
       (.I0(core_n_1517),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[43]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[47]_i_2 
       (.I0(core_n_1510),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[47]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[47]_i_3 
       (.I0(core_n_1511),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[47]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[47]_i_4 
       (.I0(core_n_1512),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[47]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[47]_i_5 
       (.I0(core_n_1513),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[47]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[51]_i_2 
       (.I0(core_n_1506),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[51]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[51]_i_3 
       (.I0(core_n_1507),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[51]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[51]_i_4 
       (.I0(core_n_1508),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[51]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[51]_i_5 
       (.I0(core_n_1509),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[51]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[55]_i_2 
       (.I0(core_n_1502),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[55]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[55]_i_3 
       (.I0(core_n_1503),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[55]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[55]_i_4 
       (.I0(core_n_1504),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[55]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[55]_i_5 
       (.I0(core_n_1505),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[55]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[59]_i_2 
       (.I0(core_n_1498),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[59]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[59]_i_3 
       (.I0(core_n_1499),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[59]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[59]_i_4 
       (.I0(core_n_1500),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[59]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[59]_i_5 
       (.I0(core_n_1501),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[59]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[63]_i_4 
       (.I0(core_n_1494),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[63]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[63]_i_5 
       (.I0(core_n_1495),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[63]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[63]_i_6 
       (.I0(core_n_1496),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[63]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAACAA)) 
    \trig_pc[63]_i_7 
       (.I0(core_n_1497),
        .I1(dcacheArb_io_requestor_1_s1_data_data[52]),
        .I2(core_n_1346),
        .I3(core_n_1345),
        .I4(core_n_1347),
        .O(\trig_pc[63]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[7]_i_2 
       (.I0(core_n_1550),
        .I1(mem_reg_pc[7]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[17]),
        .O(\trig_pc[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[7]_i_3 
       (.I0(core_n_1551),
        .I1(mem_reg_pc[6]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[16]),
        .O(\trig_pc[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[7]_i_4 
       (.I0(core_n_1552),
        .I1(mem_reg_pc[5]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[12]),
        .O(\trig_pc[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h66666F6666666066)) 
    \trig_pc[7]_i_5 
       (.I0(core_n_1553),
        .I1(mem_reg_pc[4]),
        .I2(core_n_1347),
        .I3(core_n_1345),
        .I4(core_n_1346),
        .I5(dcacheArb_io_requestor_1_s1_data_data[11]),
        .O(\trig_pc[7]_i_5_n_0 ));
  CARRY4 \trig_pc_reg[11]_i_1 
       (.CI(\trig_pc_reg[7]_i_1_n_0 ),
        .CO({\trig_pc_reg[11]_i_1_n_0 ,\trig_pc_reg[11]_i_1_n_1 ,\trig_pc_reg[11]_i_1_n_2 ,\trig_pc_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__213_n_0,core__212_n_0,core__211_n_0,core__210_n_0}),
        .O({\trig_pc_reg[11]_i_1_n_4 ,\trig_pc_reg[11]_i_1_n_5 ,\trig_pc_reg[11]_i_1_n_6 ,\trig_pc_reg[11]_i_1_n_7 }),
        .S({\trig_pc[11]_i_2_n_0 ,\trig_pc[11]_i_3_n_0 ,\trig_pc[11]_i_4_n_0 ,\trig_pc[11]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[15]_i_1 
       (.CI(\trig_pc_reg[11]_i_1_n_0 ),
        .CO({\trig_pc_reg[15]_i_1_n_0 ,\trig_pc_reg[15]_i_1_n_1 ,\trig_pc_reg[15]_i_1_n_2 ,\trig_pc_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__217_n_0,core__216_n_0,core__215_n_0,core__214_n_0}),
        .O({\trig_pc_reg[15]_i_1_n_4 ,\trig_pc_reg[15]_i_1_n_5 ,\trig_pc_reg[15]_i_1_n_6 ,\trig_pc_reg[15]_i_1_n_7 }),
        .S({\trig_pc[15]_i_2_n_0 ,\trig_pc[15]_i_3_n_0 ,\trig_pc[15]_i_4_n_0 ,\trig_pc[15]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[19]_i_1 
       (.CI(\trig_pc_reg[15]_i_1_n_0 ),
        .CO({\trig_pc_reg[19]_i_1_n_0 ,\trig_pc_reg[19]_i_1_n_1 ,\trig_pc_reg[19]_i_1_n_2 ,\trig_pc_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__221_n_0,core__220_n_0,core__219_n_0,core__218_n_0}),
        .O({\trig_pc_reg[19]_i_1_n_4 ,\trig_pc_reg[19]_i_1_n_5 ,\trig_pc_reg[19]_i_1_n_6 ,\trig_pc_reg[19]_i_1_n_7 }),
        .S({\trig_pc[19]_i_2_n_0 ,\trig_pc[19]_i_3_n_0 ,\trig_pc[19]_i_4_n_0 ,\trig_pc[19]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[23]_i_1 
       (.CI(\trig_pc_reg[19]_i_1_n_0 ),
        .CO({\trig_pc_reg[23]_i_1_n_0 ,\trig_pc_reg[23]_i_1_n_1 ,\trig_pc_reg[23]_i_1_n_2 ,\trig_pc_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__225_n_0,core__224_n_0,core__223_n_0,core__222_n_0}),
        .O({\trig_pc_reg[23]_i_1_n_4 ,\trig_pc_reg[23]_i_1_n_5 ,\trig_pc_reg[23]_i_1_n_6 ,\trig_pc_reg[23]_i_1_n_7 }),
        .S({\trig_pc[23]_i_2_n_0 ,\trig_pc[23]_i_3_n_0 ,\trig_pc[23]_i_4_n_0 ,\trig_pc[23]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[27]_i_1 
       (.CI(\trig_pc_reg[23]_i_1_n_0 ),
        .CO({\trig_pc_reg[27]_i_1_n_0 ,\trig_pc_reg[27]_i_1_n_1 ,\trig_pc_reg[27]_i_1_n_2 ,\trig_pc_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__229_n_0,core__228_n_0,core__227_n_0,core__226_n_0}),
        .O({\trig_pc_reg[27]_i_1_n_4 ,\trig_pc_reg[27]_i_1_n_5 ,\trig_pc_reg[27]_i_1_n_6 ,\trig_pc_reg[27]_i_1_n_7 }),
        .S({\trig_pc[27]_i_2_n_0 ,\trig_pc[27]_i_3_n_0 ,\trig_pc[27]_i_4_n_0 ,\trig_pc[27]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[31]_i_1 
       (.CI(\trig_pc_reg[27]_i_1_n_0 ),
        .CO({\trig_pc_reg[31]_i_1_n_0 ,\trig_pc_reg[31]_i_1_n_1 ,\trig_pc_reg[31]_i_1_n_2 ,\trig_pc_reg[31]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__233_n_0,core__232_n_0,core__231_n_0,core__230_n_0}),
        .O({\trig_pc_reg[31]_i_1_n_4 ,\trig_pc_reg[31]_i_1_n_5 ,\trig_pc_reg[31]_i_1_n_6 ,\trig_pc_reg[31]_i_1_n_7 }),
        .S({\trig_pc[31]_i_2_n_0 ,\trig_pc[31]_i_3_n_0 ,\trig_pc[31]_i_4_n_0 ,\trig_pc[31]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[35]_i_1 
       (.CI(\trig_pc_reg[31]_i_1_n_0 ),
        .CO({\trig_pc_reg[35]_i_1_n_0 ,\trig_pc_reg[35]_i_1_n_1 ,\trig_pc_reg[35]_i_1_n_2 ,\trig_pc_reg[35]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__237_n_0,core__236_n_0,core__235_n_0,core__234_n_0}),
        .O({\trig_pc_reg[35]_i_1_n_4 ,\trig_pc_reg[35]_i_1_n_5 ,\trig_pc_reg[35]_i_1_n_6 ,\trig_pc_reg[35]_i_1_n_7 }),
        .S({\trig_pc[35]_i_2_n_0 ,\trig_pc[35]_i_3_n_0 ,\trig_pc[35]_i_4_n_0 ,\trig_pc[35]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[39]_i_1 
       (.CI(\trig_pc_reg[35]_i_1_n_0 ),
        .CO({\trig_pc_reg[39]_i_1_n_0 ,\trig_pc_reg[39]_i_1_n_1 ,\trig_pc_reg[39]_i_1_n_2 ,\trig_pc_reg[39]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__241_n_0,core__240_n_0,core__239_n_0,core__238_n_0}),
        .O({\trig_pc_reg[39]_i_1_n_4 ,\trig_pc_reg[39]_i_1_n_5 ,\trig_pc_reg[39]_i_1_n_6 ,\trig_pc_reg[39]_i_1_n_7 }),
        .S({\trig_pc[39]_i_2_n_0 ,\trig_pc[39]_i_3_n_0 ,\trig_pc[39]_i_4_n_0 ,\trig_pc[39]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\trig_pc_reg[3]_i_1_n_0 ,\trig_pc_reg[3]_i_1_n_1 ,\trig_pc_reg[3]_i_1_n_2 ,\trig_pc_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__205_n_0,core__204_n_0,core__203_n_0,core__202_n_0}),
        .O({\trig_pc_reg[3]_i_1_n_4 ,\trig_pc_reg[3]_i_1_n_5 ,\trig_pc_reg[3]_i_1_n_6 ,\trig_pc_reg[3]_i_1_n_7 }),
        .S({\trig_pc[3]_i_2_n_0 ,\trig_pc[3]_i_3_n_0 ,\trig_pc[3]_i_4_n_0 ,core_rep__34_n_0}));
  CARRY4 \trig_pc_reg[43]_i_1 
       (.CI(\trig_pc_reg[39]_i_1_n_0 ),
        .CO({\trig_pc_reg[43]_i_1_n_0 ,\trig_pc_reg[43]_i_1_n_1 ,\trig_pc_reg[43]_i_1_n_2 ,\trig_pc_reg[43]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__245_n_0,core__244_n_0,core__243_n_0,core__242_n_0}),
        .O({\trig_pc_reg[43]_i_1_n_4 ,\trig_pc_reg[43]_i_1_n_5 ,\trig_pc_reg[43]_i_1_n_6 ,\trig_pc_reg[43]_i_1_n_7 }),
        .S({\trig_pc[43]_i_2_n_0 ,\trig_pc[43]_i_3_n_0 ,\trig_pc[43]_i_4_n_0 ,\trig_pc[43]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[47]_i_1 
       (.CI(\trig_pc_reg[43]_i_1_n_0 ),
        .CO({\trig_pc_reg[47]_i_1_n_0 ,\trig_pc_reg[47]_i_1_n_1 ,\trig_pc_reg[47]_i_1_n_2 ,\trig_pc_reg[47]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__249_n_0,core__248_n_0,core__247_n_0,core__246_n_0}),
        .O({\trig_pc_reg[47]_i_1_n_4 ,\trig_pc_reg[47]_i_1_n_5 ,\trig_pc_reg[47]_i_1_n_6 ,\trig_pc_reg[47]_i_1_n_7 }),
        .S({\trig_pc[47]_i_2_n_0 ,\trig_pc[47]_i_3_n_0 ,\trig_pc[47]_i_4_n_0 ,\trig_pc[47]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[51]_i_1 
       (.CI(\trig_pc_reg[47]_i_1_n_0 ),
        .CO({\trig_pc_reg[51]_i_1_n_0 ,\trig_pc_reg[51]_i_1_n_1 ,\trig_pc_reg[51]_i_1_n_2 ,\trig_pc_reg[51]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__253_n_0,core__252_n_0,core__251_n_0,core__250_n_0}),
        .O({\trig_pc_reg[51]_i_1_n_4 ,\trig_pc_reg[51]_i_1_n_5 ,\trig_pc_reg[51]_i_1_n_6 ,\trig_pc_reg[51]_i_1_n_7 }),
        .S({\trig_pc[51]_i_2_n_0 ,\trig_pc[51]_i_3_n_0 ,\trig_pc[51]_i_4_n_0 ,\trig_pc[51]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[55]_i_1 
       (.CI(\trig_pc_reg[51]_i_1_n_0 ),
        .CO({\trig_pc_reg[55]_i_1_n_0 ,\trig_pc_reg[55]_i_1_n_1 ,\trig_pc_reg[55]_i_1_n_2 ,\trig_pc_reg[55]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__257_n_0,core__256_n_0,core__255_n_0,core__254_n_0}),
        .O({\trig_pc_reg[55]_i_1_n_4 ,\trig_pc_reg[55]_i_1_n_5 ,\trig_pc_reg[55]_i_1_n_6 ,\trig_pc_reg[55]_i_1_n_7 }),
        .S({\trig_pc[55]_i_2_n_0 ,\trig_pc[55]_i_3_n_0 ,\trig_pc[55]_i_4_n_0 ,\trig_pc[55]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[59]_i_1 
       (.CI(\trig_pc_reg[55]_i_1_n_0 ),
        .CO({\trig_pc_reg[59]_i_1_n_0 ,\trig_pc_reg[59]_i_1_n_1 ,\trig_pc_reg[59]_i_1_n_2 ,\trig_pc_reg[59]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__261_n_0,core__260_n_0,core__259_n_0,core__258_n_0}),
        .O({\trig_pc_reg[59]_i_1_n_4 ,\trig_pc_reg[59]_i_1_n_5 ,\trig_pc_reg[59]_i_1_n_6 ,\trig_pc_reg[59]_i_1_n_7 }),
        .S({\trig_pc[59]_i_2_n_0 ,\trig_pc[59]_i_3_n_0 ,\trig_pc[59]_i_4_n_0 ,\trig_pc[59]_i_5_n_0 }));
  CARRY4 \trig_pc_reg[63]_i_10 
       (.CI(\trig_pc_reg[63]_i_15_n_0 ),
        .CO({\trig_pc_reg[63]_i_10_n_0 ,\trig_pc_reg[63]_i_10_n_1 ,\trig_pc_reg[63]_i_10_n_2 ,\trig_pc_reg[63]_i_10_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1481,core_n_1482,core_n_1483,core_n_1484}));
  CARRY4 \trig_pc_reg[63]_i_15 
       (.CI(\trig_pc_reg[63]_i_20_n_0 ),
        .CO({\trig_pc_reg[63]_i_15_n_0 ,\trig_pc_reg[63]_i_15_n_1 ,\trig_pc_reg[63]_i_15_n_2 ,\trig_pc_reg[63]_i_15_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1477,core_n_1478,core_n_1479,core_n_1480}));
  CARRY4 \trig_pc_reg[63]_i_2 
       (.CI(\trig_pc_reg[59]_i_1_n_0 ),
        .CO({\trig_pc_reg[63]_i_2_n_1 ,\trig_pc_reg[63]_i_2_n_2 ,\trig_pc_reg[63]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,core__264_n_0,core__263_n_0,core__262_n_0}),
        .O({\trig_pc_reg[63]_i_2_n_4 ,\trig_pc_reg[63]_i_2_n_5 ,\trig_pc_reg[63]_i_2_n_6 ,\trig_pc_reg[63]_i_2_n_7 }),
        .S({\trig_pc[63]_i_4_n_0 ,\trig_pc[63]_i_5_n_0 ,\trig_pc[63]_i_6_n_0 ,\trig_pc[63]_i_7_n_0 }));
  CARRY4 \trig_pc_reg[63]_i_20 
       (.CI(\trig_pc_reg[63]_i_25_n_0 ),
        .CO({\trig_pc_reg[63]_i_20_n_0 ,\trig_pc_reg[63]_i_20_n_1 ,\trig_pc_reg[63]_i_20_n_2 ,\trig_pc_reg[63]_i_20_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1473,core_n_1474,core_n_1475,core_n_1476}));
  CARRY4 \trig_pc_reg[63]_i_25 
       (.CI(\<const0> ),
        .CO({\trig_pc_reg[63]_i_25_n_0 ,\trig_pc_reg[63]_i_25_n_1 ,\trig_pc_reg[63]_i_25_n_2 ,\trig_pc_reg[63]_i_25_n_3 }),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1469,core_n_1470,core_n_1471,core_n_1472}));
  CARRY4 \trig_pc_reg[63]_i_3 
       (.CI(\trig_pc_reg[63]_i_8_n_0 ),
        .CO({trigB,\trig_pc_reg[63]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,core__432_n_0,core_n_1489}));
  CARRY4 \trig_pc_reg[63]_i_8 
       (.CI(\trig_pc_reg[63]_i_10_n_0 ),
        .CO({\trig_pc_reg[63]_i_8_n_0 ,\trig_pc_reg[63]_i_8_n_1 ,\trig_pc_reg[63]_i_8_n_2 ,\trig_pc_reg[63]_i_8_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1485,core_n_1486,core_n_1487,core_n_1488}));
  CARRY4 \trig_pc_reg[7]_i_1 
       (.CI(\trig_pc_reg[3]_i_1_n_0 ),
        .CO({\trig_pc_reg[7]_i_1_n_0 ,\trig_pc_reg[7]_i_1_n_1 ,\trig_pc_reg[7]_i_1_n_2 ,\trig_pc_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({core__209_n_0,core__208_n_0,core__207_n_0,core__206_n_0}),
        .O({\trig_pc_reg[7]_i_1_n_4 ,\trig_pc_reg[7]_i_1_n_5 ,\trig_pc_reg[7]_i_1_n_6 ,\trig_pc_reg[7]_i_1_n_7 }),
        .S({\trig_pc[7]_i_2_n_0 ,\trig_pc[7]_i_3_n_0 ,\trig_pc[7]_i_4_n_0 ,\trig_pc[7]_i_5_n_0 }));
  CARRY4 \trig_state_reg[1]_i_12 
       (.CI(\trig_state_reg[1]_i_17_n_0 ),
        .CO({\trig_state_reg[1]_i_12_n_0 ,\trig_state_reg[1]_i_12_n_1 ,\trig_state_reg[1]_i_12_n_2 ,\trig_state_reg[1]_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1456,core_n_1457,core_n_1458,core_n_1459}));
  CARRY4 \trig_state_reg[1]_i_17 
       (.CI(\trig_state_reg[1]_i_22_n_0 ),
        .CO({\trig_state_reg[1]_i_17_n_0 ,\trig_state_reg[1]_i_17_n_1 ,\trig_state_reg[1]_i_17_n_2 ,\trig_state_reg[1]_i_17_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1452,core_n_1453,core_n_1454,core_n_1455}));
  CARRY4 \trig_state_reg[1]_i_22 
       (.CI(\<const0> ),
        .CO({\trig_state_reg[1]_i_22_n_0 ,\trig_state_reg[1]_i_22_n_1 ,\trig_state_reg[1]_i_22_n_2 ,\trig_state_reg[1]_i_22_n_3 }),
        .CYINIT(\<const1> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1446,core_n_1447,core_n_1448,core_n_1449}));
  CARRY4 \trig_state_reg[1]_i_3 
       (.CI(\trig_state_reg[1]_i_5_n_0 ),
        .CO({trigA,\trig_state_reg[1]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({\<const0> ,\<const0> ,core__431_n_0,core_n_1468}));
  CARRY4 \trig_state_reg[1]_i_5 
       (.CI(\trig_state_reg[1]_i_7_n_0 ),
        .CO({\trig_state_reg[1]_i_5_n_0 ,\trig_state_reg[1]_i_5_n_1 ,\trig_state_reg[1]_i_5_n_2 ,\trig_state_reg[1]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1464,core_n_1465,core_n_1466,core_n_1467}));
  CARRY4 \trig_state_reg[1]_i_7 
       (.CI(\trig_state_reg[1]_i_12_n_0 ),
        .CO({\trig_state_reg[1]_i_7_n_0 ,\trig_state_reg[1]_i_7_n_1 ,\trig_state_reg[1]_i_7_n_2 ,\trig_state_reg[1]_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .S({core_n_1460,core_n_1461,core_n_1462,core_n_1463}));
endmodule 