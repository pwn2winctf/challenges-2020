module Rocket
   (req_dw_reg,
    _T_1790,
    mem_ctrl_mem,
    mem_ctrl_fp,
    wb_ctrl_mem,
    ex_ctrl_jalr,
    ex_reg_flush_pipe,
    ex_ctrl_wxd,
    ex_ctrl_div,
    mem_reg_valid,
    ex_reg_xcpt_interrupt,
    mem_reg_xcpt_interrupt,
    wb_ctrl_wxd,
    mem_ctrl_jalr,
    mem_ctrl_jal,
    mem_reg_rvc,
    mem_reg_rvc_reg_0,
    ex_reg_xcpt,
    mem_reg_xcpt,
    wb_reg_xcpt,
    wb_reg_replay,
    wb_reg_valid,
    wb_ctrl_div,
    ex_reg_valid,
    mem_ctrl_branch,
    _T_1844,
    mem_reg_sfence,
    ex_ctrl_fence_i,
    wb_ctrl_fence_i_reg_0,
    mem_reg_flush_pipe,
    \trig_pc_reg[0]_0 ,
    mem_reg_slow_bypass,
    ex_reg_rs_bypass_0_reg_0,
    _T_4899,
    \reg_mtvec_reg[20] ,
    \reg_mtvec_reg[21] ,
    \reg_mtvec_reg[22] ,
    reg_dcsr_step,
    _T_5044,
    csr_io_bp_0_control_u,
    csr_io_bp_0_control_s,
    csr_io_bp_0_control_m,
    csr_io_bp_0_control_action,
    \_T_294_reg[3] ,
    \_T_281_reg[3] ,
    csr_io_status_debug,
    reg_mstatus_spie_reg,
    reg_mstatus_mpie_reg,
    dcache_io_ptw_status_sum,
    dcache_io_ptw_status_mxr,
    reg_singleStepped,
    frontend_io_ptw_pmp_1_cfg_w,
    D,
    buf__replay,
    \ex_ctrl_sel_alu2_reg[1]_0 ,
    buf__xcpt_ae_inst,
    _T_100,
    \remainder_reg[129] ,
    \remainder_reg[129]_0 ,
    _T_216,
    \state_reg[2] ,
    Q,
    \count_reg[0] ,
    resHi_reg,
    \remainder_reg[65] ,
    \ex_reg_rs_msb_1_reg[29]_0 ,
    \remainder_reg[31] ,
    \remainder_reg[59] ,
    \s1_req_addr_reg[39] ,
    O,
    \divisor_reg[57] ,
    \remainder_reg[33] ,
    \remainder_reg[34] ,
    \remainder_reg[35] ,
    \remainder_reg[36] ,
    \remainder_reg[37] ,
    \remainder_reg[38] ,
    \remainder_reg[39] ,
    \remainder_reg[41] ,
    \remainder_reg[42] ,
    \remainder_reg[43] ,
    \remainder_reg[44] ,
    \remainder_reg[46] ,
    \remainder_reg[47] ,
    \remainder_reg[49] ,
    \remainder_reg[50] ,
    \remainder_reg[51] ,
    \remainder_reg[52] ,
    \remainder_reg[54] ,
    \remainder_reg[55] ,
    \remainder_reg[57] ,
    \remainder_reg[58] ,
    \remainder_reg[60] ,
    \remainder_reg[61] ,
    \remainder_reg[62] ,
    neg_out_reg,
    \ex_reg_rs_msb_0_reg[27]_0 ,
    \remainder_reg[63] ,
    \remainder_reg[107] ,
    \remainder_reg[111] ,
    \remainder_reg[115] ,
    \remainder_reg[119] ,
    \remainder_reg[127] ,
    \remainder_reg[127]_0 ,
    \remainder_reg[127]_1 ,
    \remainder_reg[127]_2 ,
    \remainder_reg[127]_3 ,
    \remainder_reg[123] ,
    \remainder_reg[127]_4 ,
    \remainder_reg[127]_5 ,
    \remainder_reg[129]_1 ,
    CO,
    \remainder_reg[91] ,
    \remainder_reg[95] ,
    \remainder_reg[99] ,
    \remainder_reg[103] ,
    \remainder_reg[115]_0 ,
    \remainder_reg[103]_0 ,
    \remainder_reg[103]_1 ,
    \remainder_reg[107]_0 ,
    \remainder_reg[111]_0 ,
    \remainder_reg[127]_6 ,
    \remainder_reg[115]_1 ,
    \reg_entries_0_reg[6] ,
    \reg_mtvec_reg[29] ,
    \reg_entries_0_reg[0] ,
    \reg_entries_0_reg[6]_0 ,
    \reg_mtvec_reg[29]_0 ,
    \s2_req_addr_reg[31] ,
    \reg_entries_0_reg[6]_1 ,
    \reg_mtvec_reg[29]_1 ,
    \reg_mtvec_reg[29]_2 ,
    \reg_entries_0_reg[6]_2 ,
    \reg_entries_0_reg[6]_3 ,
    \reg_entries_0_reg[6]_4 ,
    \reg_mtvec_reg[29]_3 ,
    \valid_reg[3] ,
    frontend_io_cpu_sfence_valid,
    \reg_mtvec_reg[29]_4 ,
    \reg_mtvec_reg[29]_5 ,
    \reg_mtvec_reg[29]_6 ,
    \reg_entries_1_reg[0] ,
    \reg_entries_1_reg[0]_0 ,
    \reg_entries_1_reg[0]_1 ,
    \reg_entries_1_reg[0]_2 ,
    \reg_entries_1_reg[0]_3 ,
    \reg_entries_1_reg[0]_4 ,
    \reg_entries_1_reg[0]_5 ,
    \reg_entries_1_reg[0]_6 ,
    s1_valid_reg,
    mem_reg_replay_reg_0,
    \reg_entries_1_reg[0]_7 ,
    dcache_io_ptw_resp_bits_homogeneous,
    .\s1_pc_reg[39] (_T_2177[24]),
    \reg_sbadaddr_reg[39] ,
    \reg_sscratch_reg[62] ,
    \reg_entries_1_reg[0]_8 ,
    invalidated_reg,
    SR,
    \valid_reg[3]_0 ,
    \valid_reg[3]_1 ,
    \valid_reg[3]_2 ,
    \valid_reg[3]_3 ,
    \valid_reg[1] ,
    \reg_entries_1_reg[0]_9 ,
    \reg_entries_0_reg[5] ,
    _T_1081,
    frontend_io_ptw_status_prv,
    \reg_entries_0_reg[5]_0 ,
    \reg_pmp_5_cfg_a_reg[1] ,
    \reg_entries_1_reg[0]_10 ,
    \reg_entries_0_reg[5]_1 ,
    \reg_pmp_4_cfg_a_reg[1] ,
    \reg_entries_1_reg[0]_11 ,
    \reg_entries_0_reg[5]_2 ,
    \reg_entries_0_reg[5]_3 ,
    frontend_io_ptw_pmp_7_cfg_a,
    \reg_entries_1_reg[0]_12 ,
    \reg_entries_0_reg[5]_4 ,
    frontend_io_ptw_pmp_6_cfg_a,
    \reg_entries_1_reg[0]_13 ,
    \reg_entries_0_reg[5]_5 ,
    frontend_io_ptw_pmp_2_cfg_a,
    \reg_entries_0_reg[5]_6 ,
    frontend_io_ptw_pmp_1_cfg_a,
    \reg_entries_1_reg[0]_14 ,
    \reg_entries_0_reg[5]_7 ,
    s2_valid_reg,
    frontend_io_ptw_ptbr_mode,
    bad_va,
    s2_tlb_resp_cacheable_reg,
    \reg_entries_0_reg[5]_8 ,
    \reg_entries_0_reg[5]_9 ,
    \reg_entries_0_reg[5]_10 ,
    \reg_entries_0_reg[5]_11 ,
    \reg_entries_0_reg[5]_12 ,
    \reg_entries_0_reg[5]_13 ,
    \reg_entries_0_reg[5]_14 ,
    \reg_entries_0_reg[5]_15 ,
    \reg_entries_0_reg[5]_16 ,
    \reg_entries_0_reg[5]_17 ,
    \reg_entries_0_reg[5]_18 ,
    \reg_entries_0_reg[5]_19 ,
    \reg_entries_0_reg[5]_20 ,
    \reg_entries_0_reg[5]_21 ,
    \reg_entries_0_reg[5]_22 ,
    \reg_entries_0_reg[5]_23 ,
    \reg_entries_0_reg[0]_0 ,
    p_13_in,
    \reg_entries_0_reg[5]_24 ,
    \reg_entries_0_reg[5]_25 ,
    \reg_entries_0_reg[5]_26 ,
    \reg_entries_0_reg[5]_27 ,
    \reg_entries_0_reg[5]_28 ,
    \reg_entries_0_reg[5]_29 ,
    \reg_entries_0_reg[5]_30 ,
    \reg_entries_0_reg[5]_31 ,
    \reg_entries_0_reg[5]_32 ,
    \reg_entries_0_reg[5]_33 ,
    \reg_entries_0_reg[5]_34 ,
    \reg_entries_0_reg[5]_35 ,
    \reg_entries_0_reg[5]_36 ,
    \reg_entries_0_reg[5]_37 ,
    \reg_entries_0_reg[5]_38 ,
    \reg_entries_0_reg[5]_39 ,
    \reg_entries_0_reg[5]_40 ,
    \reg_entries_0_reg[5]_41 ,
    \reg_entries_0_reg[5]_42 ,
    \reg_entries_0_reg[5]_43 ,
    \reg_entries_0_reg[5]_44 ,
    \reg_entries_0_reg[5]_45 ,
    \reg_entries_0_reg[5]_46 ,
    \reg_entries_0_reg[5]_47 ,
    \reg_entries_0_reg[0]_1 ,
    \reg_entries_0_reg[0]_2 ,
    \reg_entries_0_reg[0]_3 ,
    \reg_entries_0_reg[0]_4 ,
    \reg_entries_0_reg[0]_5 ,
    \reg_entries_0_reg[0]_6 ,
    \reg_entries_0_reg[0]_7 ,
    \ex_ctrl_sel_alu2_reg[1]_1 ,
    \ex_ctrl_sel_alu2_reg[1]_2 ,
    \ex_ctrl_sel_alu2_reg[1]_3 ,
    _T_5074,
    \_T_294_reg[0] ,
    reg_mip_seip_reg,
    \reg_pmp_7_addr_reg[29] ,
    \reg_mtvec_reg[12] ,
    \reg_sscratch_reg[59] ,
    \_T_1883_reg[1] ,
    \reg_mbadaddr_reg[12] ,
    \reg_mie_reg[7] ,
    \mem_reg_rs2_reg[7]_0 ,
    \s1_pc_reg[4] ,
    \mem_reg_rs2_reg[6]_0 ,
    \reg_sepc_reg[12] ,
    \reg_mtvec_reg[8] ,
    \reg_mepc_reg[12] ,
    reg_mip_seip_reg_0,
    \s1_pc_reg[4]_0 ,
    \reg_mtvec_reg[10] ,
    \reg_mtvec_reg[11] ,
    \reg_mtvec_reg[13] ,
    \reg_sscratch_reg[45] ,
    \r_pte_ppn_reg[19] ,
    \reg_mtvec_reg[14] ,
    \reg_mtvec_reg[15] ,
    \reg_mtvec_reg[16] ,
    \reg_mtvec_reg[17] ,
    \reg_mtvec_reg[18] ,
    \reg_mtvec_reg[19] ,
    \reg_mtvec_reg[20]_0 ,
    \reg_dpc_reg[12] ,
    \reg_mtvec_reg[21]_0 ,
    \reg_mtvec_reg[22]_0 ,
    \reg_mtvec_reg[23] ,
    \reg_mtvec_reg[24] ,
    \reg_mtvec_reg[25] ,
    \reg_mtvec_reg[26] ,
    \reg_mtvec_reg[27] ,
    \reg_mtvec_reg[28] ,
    \reg_mtvec_reg[29]_7 ,
    \reg_dscratch_reg[0] ,
    \mem_reg_rs2_reg[0]_0 ,
    \mem_reg_rs2_reg[1]_0 ,
    \reg_misa_reg[12] ,
    \mem_reg_rs2_reg[2]_0 ,
    \reg_mcause_reg[0] ,
    \mem_reg_rs2_reg[3]_0 ,
    \mem_reg_rs2_reg[4]_0 ,
    \mem_reg_rs2_reg[5]_0 ,
    csr_io_tval,
    \reg_stvec_reg[38] ,
    \reg_stvec_reg[37] ,
    \reg_stvec_reg[36] ,
    \reg_stvec_reg[35] ,
    \reg_stvec_reg[34] ,
    \reg_stvec_reg[33] ,
    \reg_stvec_reg[32] ,
    \reg_mtvec_reg[31] ,
    \reg_mtvec_reg[30] ,
    \reg_sscratch_reg[0] ,
    \reg_bp_0_control_tmatch_reg[1] ,
    \reg_sbadaddr_reg[0] ,
    \ex_cause_reg[1]_0 ,
    \reg_misa_reg[0] ,
    \reg_scause_reg[0] ,
    \reg_pmp_2_addr_reg[29] ,
    \_T_294_reg[0]_0 ,
    reg_mstatus_mie,
    reg_mstatus_mie_reg,
    \reg_sscratch_reg[45]_0 ,
    \reg_sptbr_ppn_reg[0] ,
    \_T_1883_reg[0] ,
    reg_debug_reg,
    \reg_mstatus_prv_reg[1] ,
    reg_mstatus_mpie_reg_0,
    \reg_mstatus_mpp_reg[1] ,
    \reg_mstatus_mpp_reg[0] ,
    reg_mstatus_mie_reg_0,
    \reg_dcsr_cause_reg[1] ,
    \reg_scause_reg[1] ,
    \s1_pc_reg[5] ,
    \reg_scause_reg[3] ,
    \reg_scause_reg[0]_0 ,
    \reg_dcsr_cause_reg[0] ,
    reg_wfi_reg,
    \reg_scause_reg[1]_0 ,
    reg_dcsr_prv,
    \reg_bp_0_control_tmatch_reg[1]_0 ,
    \reg_scause_reg[2] ,
    \reg_sepc_reg[26] ,
    _T_481,
    dcacheArb_io_requestor_1_req_valid,
    \s1_req_cmd_reg[4] ,
    \state_reg[1] ,
    \s1_pc_reg[1] ,
    \s1_pc_reg[39]_0 ,
    ibuf_io_inst_0_bits_xcpt0_ae_inst,
    \ex_reg_pc_reg[39]_0 ,
    \ex_ctrl_sel_alu2_reg[1]_4 ,
    ex_ctrl_mem_reg_0,
    id_reg_fence_reg_0,
    ex_ctrl_mem_reg_1,
    ex_reg_rs_bypass_1_reg_0,
    \ex_reg_rs_lsb_0_reg[0]_0 ,
    \_T_2547_reg[1]_0 ,
    ex_ctrl_mem_reg_2,
    \ex_ctrl_sel_alu2_reg[1]_5 ,
    ex_ctrl_mem_reg_3,
    ex_ctrl_mem_reg_4,
    ex_ctrl_mem_reg_5,
    _T_1829,
    \ex_reg_rs_lsb_0_reg[0]_1 ,
    \wb_reg_inst_reg[31]_0 ,
    ex_ctrl_mem_reg_6,
    \ex_reg_rs_lsb_0_reg[1]_0 ,
    _T_1406,
    _GEN_274,
    \_T_2547_reg[16]_0 ,
    ex_ctrl_mem_reg_7,
    ex_ctrl_mem_reg_8,
    ex_ctrl_mem_reg_9,
    \mem_reg_inst_reg[31]_0 ,
    \ex_reg_rs_msb_1_reg[61]_0 ,
    _T_1416,
    p_31_in,
    \ex_reg_rs_msb_1_reg[61]_1 ,
    ex_reg_rvc_reg_0,
    _T_134,
    \ex_reg_rs_msb_0_reg[10]_0 ,
    \ex_reg_rs_msb_0_reg[8]_0 ,
    \ex_reg_rs_msb_0_reg[9]_0 ,
    \ex_reg_rs_msb_0_reg[11]_0 ,
    \ex_reg_rs_msb_0_reg[12]_0 ,
    \ex_reg_rs_msb_0_reg[13]_0 ,
    \ex_reg_rs_msb_0_reg[14]_0 ,
    \ex_reg_rs_msb_0_reg[15]_0 ,
    \ex_reg_rs_msb_0_reg[16]_0 ,
    \ex_reg_rs_msb_0_reg[17]_0 ,
    \ex_reg_rs_msb_0_reg[18]_0 ,
    \ex_reg_rs_msb_0_reg[19]_0 ,
    \ex_reg_rs_msb_0_reg[20]_0 ,
    \ex_reg_rs_msb_0_reg[21]_0 ,
    \ex_reg_rs_msb_0_reg[22]_0 ,
    \ex_reg_rs_msb_0_reg[23]_0 ,
    \ex_reg_rs_msb_0_reg[24]_0 ,
    \ex_reg_rs_msb_0_reg[25]_0 ,
    \ex_reg_rs_msb_0_reg[26]_0 ,
    \ex_reg_rs_msb_0_reg[27]_1 ,
    \reg_dpc_reg[39] ,
    mem_reg_valid_reg_0,
    dcacheArb_io_requestor_1_s1_kill,
    frontend_io_cpu_req_bits_speculative,
    \wb_reg_cause_reg[0]_0 ,
    \wb_reg_cause_reg[3]_0 ,
    \ex_reg_rs_msb_1_reg[61]_2 ,
    \_T_2547_reg[31]_0 ,
    \bypass_mux_2_reg[38]_0 ,
    \mem_reg_rs2_reg[3]_1 ,
    \reg_sbadaddr_reg[30] ,
    \reg_sbadaddr_reg[30]_0 ,
    \reg_sbadaddr_reg[30]_1 ,
    \reg_sbadaddr_reg[30]_2 ,
    \lrscCount_reg[0] ,
    \lrscCount_reg[0]_0 ,
    \trig_state_reg[1]_0 ,
    \trig_state_reg[0]_0 ,
    \trig_state_reg[1]_1 ,
    \trig_state_reg[1]_2 ,
    \trig_pc_reg[0]_1 ,
    trig_pc_valid_reg_0,
    \wb_reg_pc_reg[34]_0 ,
    \bypass_mux_2_reg[35]_0 ,
    \bypass_mux_2_reg[31]_0 ,
    ex_ctrl_mem_reg_10,
    _T_1573,
    ex_ctrl_mem_reg_11,
    ex_sfence,
    mem_reg_sfence_reg_0,
    \trig_jalr_count_reg[0]_0 ,
    \a_data_reg[63] ,
    \s1_pc_reg[39]_1 ,
    \s1_pc_reg[39]_2 ,
    \s1_pc_reg[39]_3 ,
    \s1_pc_reg[39]_4 ,
    \trig_state_reg[1]_3 ,
    \trig_mem_data_reg[126]_0 ,
    \trig_state_reg[1]_4 ,
    \trig_state_reg[1]_5 ,
    \trig_state_reg[1]_6 ,
    \trig_state_reg[1]_7 ,
    \trig_state_reg[1]_8 ,
    \trig_jalr_count_reg[0]_1 ,
    \trig_jalr_count_reg[0]_2 ,
    \trig_jalr_count_reg[0]_3 ,
    \trig_jalr_count_reg[0]_4 ,
    \trig_jalr_count_reg[0]_5 ,
    \trig_jalr_count_reg[0]_6 ,
    \trig_pc_reg[0]_2 ,
    \trig_pc_reg[63]_0 ,
    \wb_reg_pc_reg[39]_0 ,
    \trig_pc_reg[0]_3 ,
    \trig_pc_reg[0]_4 ,
    \trig_pc_reg[0]_5 ,
    \trig_pc_reg[0]_6 ,
    \trig_pc_reg[0]_7 ,
    \s1_req_addr_reg[39]_0 ,
    \s1_req_addr_reg[39]_1 ,
    alu_io_in1,
    \mem_reg_pc_reg[31]_0 ,
    \ex_ctrl_sel_alu1_reg[1]_0 ,
    \ex_ctrl_sel_alu1_reg[0]_0 ,
    \remainder_reg[33]_0 ,
    \remainder_reg[34]_0 ,
    \remainder_reg[35]_0 ,
    \remainder_reg[36]_0 ,
    \remainder_reg[37]_0 ,
    \remainder_reg[38]_0 ,
    \s1_req_addr_reg[39]_2 ,
    \s1_req_addr_reg[39]_3 ,
    \reg_sbadaddr_reg[39]_0 ,
    \reg_sbadaddr_reg[39]_1 ,
    \reg_sbadaddr_reg[39]_2 ,
    \s1_pc_reg[39]_5 ,
    mem_reg_slow_bypass_reg_0,
    dcacheArb_io_requestor_1_req_bits_typ,
    alu_io_in2,
    ex_ctrl_sel_alu2,
    \mem_reg_rs2_reg[25]_0 ,
    \bypass_mux_1_reg[6]_0 ,
    \bypass_mux_1_reg[4]_0 ,
    \reg_sbadaddr_reg[30]_3 ,
    \bypass_mux_1_reg[6]_1 ,
    \bypass_mux_1_reg[0]_0 ,
    \reg_sbadaddr_reg[30]_4 ,
    \s1_req_addr_reg[3] ,
    \s1_req_addr_reg[39]_4 ,
    \reg_sbadaddr_reg[30]_5 ,
    \reg_sbadaddr_reg[30]_6 ,
    \reg_sbadaddr_reg[30]_7 ,
    \reg_sbadaddr_reg[30]_8 ,
    \reg_sbadaddr_reg[30]_9 ,
    \_T_389_reg[7] ,
    \reg_entries_1_reg[0]_15 ,
    \reg_entries_1_reg[0]_16 ,
    \reg_entries_1_reg[0]_17 ,
    \reg_entries_1_reg[0]_18 ,
    \reg_entries_1_reg[0]_19 ,
    \reg_entries_1_reg[0]_20 ,
    \reg_entries_1_reg[0]_21 ,
    \reg_entries_1_reg[0]_22 ,
    \reg_entries_1_reg[0]_23 ,
    \reg_entries_1_reg[0]_24 ,
    \reg_entries_1_reg[0]_25 ,
    \reg_entries_1_reg[0]_26 ,
    \reg_entries_1_reg[0]_27 ,
    \reg_entries_1_reg[0]_28 ,
    \reg_entries_1_reg[0]_29 ,
    \reg_entries_1_reg[0]_30 ,
    \reg_entries_1_reg[0]_31 ,
    \reg_entries_1_reg[0]_32 ,
    \reg_entries_1_reg[0]_33 ,
    \reg_entries_1_reg[0]_34 ,
    \reg_entries_1_reg[0]_35 ,
    \reg_entries_1_reg[0]_36 ,
    \reg_entries_1_reg[0]_37 ,
    \reg_entries_1_reg[0]_38 ,
    \reg_entries_1_reg[0]_39 ,
    \reg_entries_1_reg[0]_40 ,
    \reg_entries_1_reg[0]_41 ,
    \reg_entries_1_reg[0]_42 ,
    \reg_entries_1_reg[0]_43 ,
    \reg_entries_1_reg[0]_44 ,
    \reg_entries_1_reg[0]_45 ,
    \reg_entries_1_reg[0]_46 ,
    \reg_entries_1_reg[0]_47 ,
    \reg_entries_0_reg[6]_5 ,
    \reg_entries_0_reg[4] ,
    \reg_entries_0_reg[6]_6 ,
    _T_4068_ae_ld_reg,
    _T_4068_pf_ld_reg,
    \valid_reg[0] ,
    \r_refill_waddr_reg[0] ,
    \_T_973_reg[1] ,
    \reg_entries_0_reg[6]_7 ,
    \reg_entries_0_reg[4]_0 ,
    \reg_entries_0_reg[4]_1 ,
    \reg_entries_0_reg[4]_2 ,
    \reg_entries_0_reg[6]_8 ,
    \reg_entries_0_reg[6]_9 ,
    \reg_entries_0_reg[6]_10 ,
    \reg_entries_0_reg[6]_11 ,
    \reg_entries_0_reg[6]_12 ,
    \reg_entries_0_reg[6]_13 ,
    \reg_entries_0_reg[6]_14 ,
    \reg_entries_0_reg[6]_15 ,
    \reg_entries_0_reg[6]_16 ,
    \reg_entries_0_reg[6]_17 ,
    \reg_entries_0_reg[4]_3 ,
    \reg_entries_0_reg[4]_4 ,
    \reg_entries_0_reg[6]_18 ,
    \reg_entries_0_reg[6]_19 ,
    \reg_entries_0_reg[6]_20 ,
    \reg_entries_0_reg[6]_21 ,
    \reg_entries_0_reg[6]_22 ,
    \reg_entries_0_reg[6]_23 ,
    \reg_entries_0_reg[6]_24 ,
    \reg_entries_0_reg[6]_25 ,
    \reg_entries_0_reg[6]_26 ,
    \reg_entries_0_reg[4]_5 ,
    \reg_entries_0_reg[4]_6 ,
    \reg_entries_0_reg[4]_7 ,
    \reg_entries_0_reg[4]_8 ,
    \reg_entries_0_reg[4]_9 ,
    \reg_entries_0_reg[6]_27 ,
    \reg_entries_0_reg[6]_28 ,
    \reg_entries_0_reg[6]_29 ,
    \reg_entries_0_reg[6]_30 ,
    \reg_entries_0_reg[6]_31 ,
    \reg_entries_0_reg[6]_32 ,
    \reg_entries_0_reg[6]_33 ,
    \reg_entries_0_reg[6]_34 ,
    \reg_entries_0_reg[6]_35 ,
    \reg_entries_0_reg[6]_36 ,
    \reg_entries_0_reg[4]_10 ,
    \reg_entries_0_reg[4]_11 ,
    \reg_entries_0_reg[4]_12 ,
    \reg_entries_0_reg[6]_37 ,
    \reg_entries_0_reg[6]_38 ,
    \reg_entries_0_reg[6]_39 ,
    \reg_entries_0_reg[4]_13 ,
    \reg_entries_0_reg[6]_40 ,
    \reg_entries_0_reg[6]_41 ,
    \reg_entries_0_reg[4]_14 ,
    \reg_entries_0_reg[4]_15 ,
    \reg_entries_0_reg[4]_16 ,
    \reg_entries_0_reg[6]_42 ,
    \reg_entries_0_reg[6]_43 ,
    \reg_entries_0_reg[6]_44 ,
    \reg_entries_0_reg[6]_45 ,
    \reg_entries_0_reg[6]_46 ,
    \reg_entries_0_reg[6]_47 ,
    \reg_entries_0_reg[6]_48 ,
    \reg_entries_0_reg[6]_49 ,
    \reg_entries_0_reg[6]_50 ,
    \reg_entries_0_reg[4]_17 ,
    \reg_entries_0_reg[6]_51 ,
    \reg_entries_0_reg[6]_52 ,
    \reg_entries_0_reg[6]_53 ,
    \reg_entries_0_reg[6]_54 ,
    \reg_entries_0_reg[6]_55 ,
    \reg_entries_0_reg[4]_18 ,
    \reg_entries_0_reg[6]_56 ,
    \reg_entries_0_reg[6]_57 ,
    \reg_entries_0_reg[4]_19 ,
    \reg_entries_0_reg[4]_20 ,
    \reg_entries_0_reg[4]_21 ,
    \reg_entries_0_reg[4]_22 ,
    \reg_entries_0_reg[4]_23 ,
    \reg_entries_0_reg[4]_24 ,
    \reg_entries_0_reg[4]_25 ,
    _T_4068_pf_ld_reg_0,
    _T_4068_pf_st_reg,
    _T_4068_pf_ld_reg_1,
    _T_4068_pf_ld_reg_2,
    _T_4068_pf_st_reg_0,
    _T_4068_pf_ld_reg_3,
    _T_4068_pf_st_reg_1,
    \ex_reg_inst_reg[11]_0 ,
    \ex_cause_reg[1]_1 ,
    \ex_cause_reg[1]_2 ,
    \ex_cause_reg[1]_3 ,
    \ex_cause_reg[1]_4 ,
    \ex_cause_reg[1]_5 ,
    \ex_cause_reg[1]_6 ,
    \ex_cause_reg[1]_7 ,
    \ex_cause_reg[1]_8 ,
    \ex_cause_reg[1]_9 ,
    \ex_cause_reg[1]_10 ,
    \ex_cause_reg[1]_11 ,
    \ex_cause_reg[1]_12 ,
    \ex_cause_reg[1]_13 ,
    \ex_cause_reg[1]_14 ,
    \wb_reg_cause_reg[0]_1 ,
    \wb_reg_cause_reg[0]_2 ,
    \wb_reg_cause_reg[0]_3 ,
    \wb_reg_cause_reg[0]_4 ,
    \wb_reg_cause_reg[0]_5 ,
    \wb_reg_cause_reg[0]_6 ,
    \wb_reg_cause_reg[0]_7 ,
    \wb_reg_cause_reg[0]_8 ,
    \wb_reg_cause_reg[0]_9 ,
    \wb_reg_cause_reg[0]_10 ,
    \wb_reg_cause_reg[0]_11 ,
    \wb_reg_cause_reg[0]_12 ,
    \wb_reg_cause_reg[0]_13 ,
    \wb_reg_cause_reg[0]_14 ,
    _T_217,
    \bypass_mux_1_reg[32]_0 ,
    \bypass_mux_1_reg[33]_0 ,
    \bypass_mux_1_reg[34]_0 ,
    \bypass_mux_1_reg[35]_0 ,
    \bypass_mux_1_reg[36]_0 ,
    \bypass_mux_1_reg[37]_0 ,
    \bypass_mux_1_reg[38]_0 ,
    \bypass_mux_1_reg[39]_0 ,
    \bypass_mux_1_reg[40]_0 ,
    \bypass_mux_1_reg[41]_0 ,
    \bypass_mux_1_reg[42]_0 ,
    \bypass_mux_1_reg[43]_0 ,
    \bypass_mux_1_reg[44]_0 ,
    \bypass_mux_1_reg[45]_0 ,
    \bypass_mux_1_reg[46]_0 ,
    \bypass_mux_1_reg[47]_0 ,
    \bypass_mux_1_reg[60]_0 ,
    \bypass_mux_1_reg[61]_0 ,
    \bypass_mux_1_reg[62]_0 ,
    \bypass_mux_1_reg[63]_0 ,
    \bypass_mux_1_reg[48]_0 ,
    \bypass_mux_1_reg[49]_0 ,
    \bypass_mux_1_reg[50]_0 ,
    \bypass_mux_1_reg[51]_0 ,
    \bypass_mux_1_reg[52]_0 ,
    \bypass_mux_1_reg[53]_0 ,
    \bypass_mux_1_reg[54]_0 ,
    \bypass_mux_1_reg[55]_0 ,
    \bypass_mux_1_reg[56]_0 ,
    \bypass_mux_1_reg[57]_0 ,
    \bypass_mux_1_reg[58]_0 ,
    \bypass_mux_1_reg[59]_0 ,
    \bypass_mux_1_reg[1]_0 ,
    shamt,
    \bypass_mux_1_reg[62]_1 ,
    \bypass_mux_1_reg[61]_1 ,
    \bypass_mux_1_reg[60]_1 ,
    \bypass_mux_1_reg[59]_1 ,
    \bypass_mux_1_reg[58]_1 ,
    \bypass_mux_1_reg[57]_1 ,
    \bypass_mux_1_reg[56]_1 ,
    \bypass_mux_1_reg[55]_1 ,
    \bypass_mux_1_reg[54]_1 ,
    \bypass_mux_1_reg[53]_1 ,
    \bypass_mux_1_reg[52]_1 ,
    \bypass_mux_1_reg[51]_1 ,
    \bypass_mux_1_reg[50]_1 ,
    \bypass_mux_1_reg[49]_1 ,
    \bypass_mux_1_reg[48]_1 ,
    \bypass_mux_1_reg[48]_2 ,
    \bypass_mux_1_reg[47]_1 ,
    \bypass_mux_1_reg[47]_2 ,
    _T_121,
    \bypass_mux_1_reg[46]_1 ,
    \bypass_mux_1_reg[46]_2 ,
    \bypass_mux_1_reg[45]_1 ,
    \bypass_mux_1_reg[45]_2 ,
    \bypass_mux_1_reg[44]_1 ,
    \bypass_mux_1_reg[44]_2 ,
    \bypass_mux_1_reg[43]_1 ,
    \bypass_mux_1_reg[43]_2 ,
    \bypass_mux_1_reg[42]_1 ,
    \bypass_mux_1_reg[42]_2 ,
    \bypass_mux_1_reg[41]_1 ,
    \bypass_mux_1_reg[41]_2 ,
    \bypass_mux_1_reg[40]_1 ,
    \bypass_mux_1_reg[40]_2 ,
    \bypass_mux_1_reg[39]_1 ,
    \bypass_mux_1_reg[39]_2 ,
    \bypass_mux_1_reg[38]_1 ,
    \bypass_mux_1_reg[38]_2 ,
    \bypass_mux_1_reg[37]_1 ,
    \bypass_mux_1_reg[37]_2 ,
    \bypass_mux_1_reg[36]_1 ,
    \bypass_mux_1_reg[35]_1 ,
    \bypass_mux_1_reg[35]_2 ,
    \bypass_mux_1_reg[34]_1 ,
    \bypass_mux_1_reg[34]_2 ,
    \bypass_mux_1_reg[33]_1 ,
    \bypass_mux_1_reg[29]_0 ,
    \bypass_mux_1_reg[33]_2 ,
    \bypass_mux_1_reg[35]_3 ,
    \bypass_mux_1_reg[29]_1 ,
    \bypass_mux_1_reg[34]_3 ,
    \bypass_mux_1_reg[34]_4 ,
    \bypass_mux_1_reg[33]_3 ,
    \bypass_mux_1_reg[33]_4 ,
    \bypass_mux_1_reg[29]_2 ,
    \bypass_mux_1_reg[29]_3 ,
    \bypass_mux_1_reg[29]_4 ,
    \bypass_mux_1_reg[23]_0 ,
    \bypass_mux_1_reg[22]_0 ,
    \bypass_mux_1_reg[21]_0 ,
    \bypass_mux_1_reg[20]_0 ,
    \bypass_mux_1_reg[19]_0 ,
    \bypass_mux_1_reg[18]_0 ,
    \bypass_mux_1_reg[17]_0 ,
    \bypass_mux_1_reg[50]_2 ,
    \bypass_mux_1_reg[51]_2 ,
    \bypass_mux_1_reg[52]_2 ,
    \bypass_mux_1_reg[53]_2 ,
    \bypass_mux_1_reg[54]_2 ,
    \bypass_mux_1_reg[55]_2 ,
    \bypass_mux_1_reg[56]_2 ,
    \bypass_mux_1_reg[57]_2 ,
    \bypass_mux_1_reg[58]_2 ,
    \bypass_mux_1_reg[59]_2 ,
    \bypass_mux_1_reg[3]_0 ,
    \bypass_mux_1_reg[2]_0 ,
    \bypass_mux_1_reg[1]_1 ,
    \bypass_mux_1_reg[1]_2 ,
    mem_br_taken__reg_0,
    \bypass_mux_1_reg[48]_3 ,
    \bypass_mux_1_reg[49]_2 ,
    \bypass_mux_1_reg[50]_3 ,
    \bypass_mux_1_reg[51]_3 ,
    \bypass_mux_1_reg[52]_3 ,
    \bypass_mux_1_reg[53]_3 ,
    \bypass_mux_1_reg[54]_3 ,
    \bypass_mux_1_reg[55]_3 ,
    \bypass_mux_1_reg[56]_3 ,
    \bypass_mux_1_reg[57]_3 ,
    \bypass_mux_1_reg[58]_3 ,
    \bypass_mux_1_reg[59]_3 ,
    host_clk,
    id_ctrl_mem,
    \buf__data_reg[1] ,
    _T_1821,
    id_ctrl_wxd,
    \buf__data_reg[1]_0 ,
    id_ctrl_jal,
    mem_reg_xcpt0,
    \buf__data_reg[1]_1 ,
    id_ctrl_rxs2,
    id_ctrl_fence_i,
    ex_ctrl_div_reg_0,
    mem_reg_flush_pipe_reg_0,
    mem_reg_sfence_reg_1,
    ex_reg_rvc_reg_1,
    target_reset,
    trig_pc_valid_reg_1,
    mem_ctrl_fence_i_reg_0,
    ex_ctrl_alu_dw_reg_0,
    mem_reg_slow_bypass_reg_1,
    ex_reg_rs_bypass_0_reg_1,
    reg_debug_reg_0,
    tile_auto_int_sync_xing_sinklzy_in_2_sync_0,
    sys_reset_reg,
    reg_debug_reg_1,
    \ex_ctrl_csr_reg[2]_0 ,
    \ex_ctrl_csr_reg[1]_0 ,
    \ex_ctrl_csr_reg[0]_0 ,
    buf__pc,
    frontend_io_cpu_resp_bits_replay,
    frontend_io_cpu_resp_bits_xcpt_pf_inst,
    frontend_io_cpu_resp_bits_xcpt_ae_inst,
    nBufValid_reg,
    \state_reg[1]_0 ,
    doUncachedResp_reg,
    \bypass_mux_2_reg[9]_0 ,
    \state_reg[0] ,
    S,
    \remainder_reg[71] ,
    \remainder_reg[75] ,
    \remainder_reg[79] ,
    \remainder_reg[83] ,
    \remainder_reg[87] ,
    \remainder_reg[91]_0 ,
    \remainder_reg[95]_0 ,
    \remainder_reg[99]_0 ,
    \remainder_reg[103]_2 ,
    \remainder_reg[107]_1 ,
    \remainder_reg[111]_1 ,
    \remainder_reg[115]_2 ,
    \remainder_reg[119]_0 ,
    \remainder_reg[123]_0 ,
    \remainder_reg[127]_7 ,
    \remainder_reg[128] ,
    \divisor_reg[35] ,
    \divisor_reg[52] ,
    \remainder_reg[64] ,
    \remainder_reg[64]_0 ,
    \remainder_reg[64]_1 ,
    \remainder_reg[64]_2 ,
    \divisor_reg[1] ,
    \divisor_reg[18] ,
    \divisor_reg[15] ,
    \divisor_reg[15]_0 ,
    \divisor_reg[15]_1 ,
    \divisor_reg[15]_2 ,
    DI,
    \divisor_reg[15]_3 ,
    \divisor_reg[15]_4 ,
    \divisor_reg[15]_5 ,
    \divisor_reg[15]_6 ,
    \divisor_reg[15]_7 ,
    \divisor_reg[15]_8 ,
    \divisor_reg[32] ,
    \remainder_reg[64]_3 ,
    \remainder_reg[64]_4 ,
    \remainder_reg[64]_5 ,
    \remainder_reg[64]_6 ,
    \divisor_reg[51] ,
    \divisor_reg[32]_0 ,
    \divisor_reg[32]_1 ,
    \remainder_reg[64]_7 ,
    \remainder_reg[64]_8 ,
    \remainder_reg[64]_9 ,
    \reg_entries_4_reg[61] ,
    \s1_req_addr_reg[31] ,
    dcache_io_ptw_resp_valid,
    \r_pte_ppn_reg[19]_0 ,
    s1_req_phys_reg,
    \reg_pmp_7_cfg_a_reg[0] ,
    s2_replay,
    \r_pte_ppn_reg[7] ,
    \r_pte_ppn_reg[7]_0 ,
    \r_pte_ppn_reg[7]_1 ,
    \r_pte_ppn_reg[7]_2 ,
    \r_pte_ppn_reg[7]_3 ,
    \r_pte_ppn_reg[7]_4 ,
    \r_pte_ppn_reg[7]_5 ,
    \r_pte_ppn_reg[7]_6 ,
    io_mask,
    dcache_io_ptw_resp_bits_ae,
    \s1_req_typ_reg[1] ,
    \r_pte_ppn_reg[5] ,
    _T_200__0,
    \s1_pc_reg[39]_6 ,
    dcacheArb_io_requestor_1_s2_nack,
    invalidated,
    refill_valid,
    p_2_in,
    _T_1432,
    \valid_reg[3]_4 ,
    \reg_entries_3_reg[11] ,
    \r_refill_waddr_reg[1] ,
    \s1_pc_reg[31] ,
    resp_valid_1_reg,
    \reg_pmp_0_addr_reg[28] ,
    _T_726,
    \reg_pmp_5_addr_reg[28] ,
    \reg_pmp_4_addr_reg[28] ,
    \reg_pmp_3_addr_reg[28] ,
    \reg_pmp_2_addr_reg[28] ,
    \reg_pmp_7_addr_reg[28] ,
    \reg_pmp_6_addr_reg[28] ,
    \reg_pmp_1_addr_reg[28] ,
    hitsVec_4,
    _T_382,
    \reg_pmp_0_addr_reg[29] ,
    \reg_pmp_1_addr_reg[29] ,
    \reg_pmp_2_addr_reg[29]_0 ,
    \reg_pmp_6_addr_reg[29] ,
    \reg_pmp_7_addr_reg[29]_0 ,
    \reg_pmp_3_addr_reg[29] ,
    \reg_pmp_4_addr_reg[29] ,
    \reg_pmp_5_addr_reg[29] ,
    _T_382__0,
    \s1_pc_reg[26] ,
    \reg_pmp_5_addr_reg[17] ,
    \reg_pmp_4_addr_reg[17] ,
    \reg_pmp_3_addr_reg[17] ,
    \reg_pmp_7_addr_reg[17] ,
    \reg_pmp_6_addr_reg[17] ,
    \reg_pmp_2_addr_reg[17] ,
    \reg_pmp_1_addr_reg[17] ,
    \reg_pmp_0_addr_reg[17] ,
    _T_480,
    \reg_pmp_5_addr_reg[19] ,
    \reg_pmp_4_addr_reg[19] ,
    \reg_pmp_3_addr_reg[19] ,
    \reg_pmp_7_addr_reg[19] ,
    \reg_pmp_6_addr_reg[19] ,
    \reg_pmp_2_addr_reg[19] ,
    \reg_pmp_1_addr_reg[19] ,
    \reg_pmp_0_addr_reg[19] ,
    \reg_pmp_5_addr_reg[13] ,
    \reg_pmp_4_addr_reg[13] ,
    \reg_pmp_3_addr_reg[13] ,
    \reg_pmp_7_addr_reg[13] ,
    \reg_pmp_6_addr_reg[13] ,
    \reg_pmp_2_addr_reg[13] ,
    \reg_pmp_1_addr_reg[13] ,
    \reg_pmp_0_addr_reg[13] ,
    nBufValid_reg_0,
    nBufValid_reg_1,
    frontend_io_cpu_resp_bits_data,
    ibuf_io_inst_0_bits_raw,
    \wb_reg_inst_reg[21]_0 ,
    \wb_reg_cause_reg[63]_0 ,
    \wb_reg_inst_reg[21]_1 ,
    \wb_reg_inst_reg[22]_0 ,
    \wb_reg_inst_reg[21]_2 ,
    \wb_reg_inst_reg[21]_3 ,
    wb_reg_replay_reg_0,
    \wb_ctrl_csr_reg[2]_0 ,
    \wb_reg_inst_reg[29]_0 ,
    tile_auto_int_sync_xing_sinklzy_in_0_sync_0,
    \wb_reg_inst_reg[21]_4 ,
    \wb_reg_inst_reg[21]_5 ,
    \reg_pmp_5_addr_reg[20] ,
    \wb_reg_inst_reg[30]_0 ,
    \wb_reg_inst_reg[30]_1 ,
    \reg_mstatus_prv_reg[1]_0 ,
    tile_auto_int_sync_xing_sinklzy_in_0_sync_1,
    tile_auto_int_sync_xing_sinklzy_in_1_sync_0,
    \wb_reg_inst_reg[29]_1 ,
    reg_debug_reg_2,
    \wb_reg_inst_reg[22]_1 ,
    \wb_reg_cause_reg[2]_0 ,
    \wb_ctrl_csr_reg[0]_0 ,
    dcache_io_cpu_invalidate_lr,
    \wb_reg_inst_reg[26]_0 ,
    \reg_mstatus_prv_reg[1]_1 ,
    wb_reg_replay_reg_1,
    \_T_294_reg[0]_1 ,
    \_T_281_reg[0] ,
    q_reg,
    \state_reg[0]_0 ,
    \state_reg[1]_1 ,
    \state_reg[0]_1 ,
    \s2_pc_reg[1] ,
    frontend_io_cpu_resp_bits_pc,
    \elts_0_pc_reg[39] ,
    nBufValid_reg_2,
    frontend_io_cpu_resp_valid,
    buf__xcpt_pf_inst_reg,
    reg_mstatus_tvm_reg,
    \s2_req_tag_reg[5] ,
    \wb_reg_inst_reg[7]_0 ,
    \buf__data_reg[3] ,
    dcacheArb_io_requestor_1_ordered,
    \buf__data_reg[2] ,
    nBufValid_reg_3,
    \buf__data_reg[4] ,
    nBufValid_reg_4,
    ibuf_io_inst_0_bits_inst_rs2,
    \buf__data_reg[3]_0 ,
    ibuf_io_inst_0_bits_inst_rs1,
    \_T_2547_reg[16]_1 ,
    nBufValid_reg_5,
    \ex_reg_inst_reg[10]_0 ,
    \wb_reg_inst_reg[7]_1 ,
    \state_reg[0]_2 ,
    \buf__data_reg[12] ,
    _T_1005,
    \mem_reg_inst_reg[11]_0 ,
    ibuf_io_inst_0_bits_inst_rd,
    \s2_req_typ_reg[0] ,
    \req_tag_reg[4] ,
    ex_ctrl_wxd_reg_0,
    reg_bp_0_control_action_reg,
    buf__xcpt_pf_inst_reg_0,
    \s2_req_cmd_reg[1] ,
    dcacheArb_io_requestor_1_resp_bits_data,
    \reg_mtvec_reg[4] ,
    wb_reg_valid_reg_0,
    dcacheArb_io_requestor_1_replay_next,
    mem_reg_sfence_reg_2,
    dcacheArb_io_requestor_1_resp_valid,
    dcacheArb_io_requestor_1_req_ready,
    wb_reg_replay_reg_2,
    \s2_req_tag_reg[5]_0 ,
    \s2_req_tag_reg[6] ,
    dcacheArb_io_requestor_1_resp_bits_replay,
    \req_tag_reg[0] ,
    \s2_req_tag_reg[6]_0 ,
    \wb_reg_inst_reg[9]_0 ,
    \req_tag_reg[1] ,
    \wb_reg_inst_reg[9]_1 ,
    \req_tag_reg[1]_0 ,
    \wb_reg_inst_reg[9]_2 ,
    \req_tag_reg[1]_1 ,
    \req_tag_reg[0]_0 ,
    \req_tag_reg[1]_2 ,
    \req_tag_reg[1]_3 ,
    \req_tag_reg[1]_4 ,
    \wb_reg_inst_reg[9]_3 ,
    p_0_in,
    dcacheArb_io_requestor_1_s2_xcpt_ma_st,
    wb_ctrl_mem_reg_0,
    dcacheArb_io_requestor_1_s2_xcpt_pf_st,
    dcacheArb_io_requestor_1_s2_xcpt_pf_ld,
    dcacheArb_io_requestor_1_s2_xcpt_ma_ld,
    \bypass_mux_2_reg[63]_0 ,
    \bypass_mux_2_reg[63]_1 ,
    \trig_mem_data_reg[127]_0 ,
    \trig_mem_data_reg[63]_0 ,
    trig_pc_valid_reg_2,
    \bypass_mux_1_reg[63]_1 ,
    \bypass_mux_1_reg[63]_2 ,
    \trig_state_reg[0]_1 ,
    \trig_pc_reg[63]_1 ,
    dcacheArb_io_requestor_1_resp_bits_data_word_bypass,
    \ex_ctrl_mem_type_reg[0]_0 ,
    \ex_ctrl_sel_imm_reg[1]_0 ,
    \wb_reg_cause_reg[63]_1 ,
    \wb_reg_cause_reg[63]_2 ,
    \wb_reg_cause_reg[63]_3 ,
    \wb_reg_cause_reg[63]_4 ,
    \wb_reg_cause_reg[63]_5 ,
    \wb_reg_cause_reg[63]_6 ,
    \ex_ctrl_sel_imm_reg[1]_1 ,
    \reg_pmp_5_cfg_a_reg[1]_0 ,
    \count_reg[1] ,
    \r_pte_ppn_reg[3] ,
    \r_pte_ppn_reg[5]_0 ,
    \r_pte_ppn_reg[16] ,
    \count_reg[1]_0 ,
    \r_pte_ppn_reg[3]_0 ,
    \r_pte_ppn_reg[5]_1 ,
    \r_pte_ppn_reg[16]_0 ,
    \r_pte_ppn_reg[3]_1 ,
    \r_pte_ppn_reg[5]_2 ,
    \r_pte_ppn_reg[16]_1 ,
    \r_pte_ppn_reg[3]_2 ,
    \r_pte_ppn_reg[5]_3 ,
    \r_pte_ppn_reg[16]_2 ,
    _T_1156,
    \r_pte_ppn_reg[3]_3 ,
    \r_pte_ppn_reg[5]_4 ,
    \r_pte_ppn_reg[16]_3 ,
    _T_931,
    \reg_pmp_0_addr_reg[28]_0 ,
    \r_pte_ppn_reg[3]_4 ,
    \r_pte_ppn_reg[5]_5 ,
    \r_pte_ppn_reg[16]_4 ,
    \count_reg[1]_1 ,
    \r_pte_ppn_reg[3]_5 ,
    \r_pte_ppn_reg[5]_6 ,
    \r_pte_ppn_reg[16]_5 ,
    \count_reg[1]_2 ,
    \r_pte_ppn_reg[3]_6 ,
    \r_pte_ppn_reg[5]_7 ,
    \r_pte_ppn_reg[16]_6 ,
    dcache_io_ptw_resp_bits_level,
    \reg_pmp_5_addr_reg[28]_0 ,
    \reg_pmp_6_addr_reg[28]_0 ,
    \reg_pmp_1_addr_reg[28]_0 ,
    \reg_pmp_2_addr_reg[28]_0 ,
    \reg_pmp_7_addr_reg[28]_0 ,
    \reg_pmp_4_addr_reg[28]_0 ,
    \reg_pmp_3_addr_reg[28]_0 ,
    s1_req_phys_reg_0,
    \reg_entries_4_reg[61]_0 ,
    \valid_reg[4] ,
    \reg_entries_0_reg[10] ,
    \valid_reg[2] ,
    \valid_reg[0]_0 ,
    \valid_reg[1]_0 ,
    \reg_pmp_1_cfg_a_reg[0] ,
    \reg_pmp_2_cfg_a_reg[0] ,
    resp_valid_0_reg,
    reg_pmp_1_cfg_w_reg,
    \s1_req_addr_reg[2] ,
    \s1_req_typ_reg[0] ,
    \s1_req_typ_reg[0]_0 ,
    tlb_io_req_bits_sfence_bits_rs2,
    \reg_pmp_1_addr_reg[29]_0 ,
    \s1_req_addr_reg[2]_0 ,
    \r_pte_ppn_reg[11] ,
    _T_382_0,
    \r_pte_ppn_reg[16]_7 ,
    \reg_pmp_3_addr_reg[29]_0 ,
    \reg_pmp_2_addr_reg[0] ,
    \reg_pmp_2_addr_reg[29]_1 ,
    \s1_req_typ_reg[0]_1 ,
    \s1_req_typ_reg[0]_2 ,
    \reg_pmp_4_addr_reg[14] ,
    \reg_pmp_4_addr_reg[0] ,
    \reg_pmp_5_addr_reg[29]_0 ,
    \s1_req_addr_reg[2]_1 ,
    \s1_req_typ_reg[0]_3 ,
    \reg_pmp_4_addr_reg[29]_0 ,
    \reg_pmp_3_addr_reg[23] ,
    \reg_pmp_3_addr_reg[29]_1 ,
    \r_pte_ppn_reg[15] ,
    \reg_pmp_6_addr_reg[29]_0 ,
    \s1_req_addr_reg[2]_2 ,
    \reg_pmp_0_addr_reg[29]_0 ,
    \reg_pmp_0_addr_reg[23] ,
    \r_pte_ppn_reg[6] ,
    \reg_pmp_7_addr_reg[29]_1 ,
    \r_pte_ppn_reg[10] ,
    \r_pte_ppn_reg[3]_7 ,
    \reg_pmp_7_addr_reg[23] ,
    \reg_pmp_7_addr_reg[29]_2 ,
    \r_pte_ppn_reg[2] ,
    \r_pte_ppn_reg[14] ,
    \r_pte_ppn_reg[7]_7 ,
    \r_pte_ppn_reg[13] ,
    \r_pte_ppn_reg[0] ,
    \r_pte_ppn_reg[8] ,
    \r_pte_ppn_reg[4] ,
    \r_pte_ppn_reg[1] ,
    \r_pte_ppn_reg[17] ,
    \r_pte_ppn_reg[18] ,
    _T_1701,
    \reg_pmp_7_addr_reg[17]_0 ,
    \r_pte_ppn_reg[9] ,
    \reg_pmp_3_addr_reg[18] ,
    \r_pte_ppn_reg[12] ,
    \reg_entries_2_reg[12] ,
    \reg_entries_1_reg[12] ,
    \reg_entries_3_reg[12] ,
    \remainder_reg[62]_0 ,
    sys_reset_reg_0,
    ADDRA,
    nBufValid_reg_6,
    _T_909,
    _T_1142,
    _T_877,
    _T_889,
    _T_1031,
    \buf__data_reg[3]_1 ,
    ex_ctrl_alu_dw_reg_1,
    ex_ctrl_alu_dw_reg_2,
    ex_ctrl_alu_dw_reg_3,
    ex_ctrl_alu_dw_reg_4,
    ex_ctrl_alu_dw_reg_5,
    ex_ctrl_alu_dw_reg_6,
    ex_ctrl_alu_dw_reg_7,
    ex_ctrl_alu_dw_reg_8,
    ex_ctrl_alu_dw_reg_9,
    ex_ctrl_alu_dw_reg_10,
    ex_ctrl_alu_dw_reg_11,
    ex_ctrl_alu_dw_reg_12,
    ex_ctrl_alu_dw_reg_13,
    ex_ctrl_alu_dw_reg_14,
    ex_ctrl_alu_dw_reg_15,
    ex_ctrl_alu_dw_reg_16,
    ex_ctrl_alu_dw_reg_17,
    ex_ctrl_alu_dw_reg_18,
    ex_ctrl_alu_dw_reg_19,
    ex_ctrl_alu_dw_reg_20,
    ex_ctrl_alu_dw_reg_21,
    ex_ctrl_alu_dw_reg_22,
    ex_ctrl_alu_dw_reg_23,
    ex_ctrl_alu_dw_reg_24,
    ex_ctrl_alu_dw_reg_25,
    ex_ctrl_alu_dw_reg_26,
    ex_ctrl_alu_dw_reg_27,
    ex_ctrl_alu_dw_reg_28,
    ex_ctrl_alu_dw_reg_29,
    ex_ctrl_alu_dw_reg_30,
    ex_ctrl_alu_dw_reg_31,
    ex_ctrl_alu_dw_reg_32,
    \buf__data_reg[1]_2 ,
    E,
    \buf__data_reg[3]_2 ,
    nBufValid_reg_7,
    ex_ctrl_wxd_reg_1,
    \mem_reg_inst_reg[9]_0 ,
    out,
    mem_ctrl_branch_reg_0,
    \buf__data_reg[1]_3 ,
    \mem_reg_inst_reg[9]_1 ,
    \bypass_mux_2_reg[63]_2 ,
    \buf__data_reg[3]_3 ,
    mem_reg_xcpt_interrupt_reg_0,
    nBufValid_reg_8,
    buf__xcpt_pf_inst_reg_1,
    \buf__data_reg[4]_0 ,
    elts_0_xcpt_ae_inst_reg,
    buf__xcpt_pf_inst_reg_2,
    \reg_misa_reg[12]_0 ,
    id_ctrl_sel_alu1,
    sys_reset_reg_1,
    sys_reset_reg_2,
    \wb_ctrl_csr_reg[0]_1 ,
    \wb_reg_pc_reg[39]_1 ,
    \wb_ctrl_csr_reg[0]_2 ,
    \wb_ctrl_csr_reg[0]_3 ,
    \wb_ctrl_csr_reg[0]_4 ,
    \wb_ctrl_csr_reg[0]_5 ,
    \wb_ctrl_csr_reg[0]_6 ,
    \wb_reg_pc_reg[39]_2 ,
    \wb_ctrl_csr_reg[0]_7 ,
    \wb_ctrl_csr_reg[0]_8 ,
    \wb_ctrl_csr_reg[0]_9 ,
    \wb_reg_pc_reg[39]_3 ,
    \wb_ctrl_csr_reg[0]_10 ,
    nBufValid_reg_9,
    \elts_0_data_reg[15] ,
    \reg_bp_0_address_reg[3] ,
    \reg_bp_0_address_reg[36] ,
    \elts_0_pc_reg[38] ,
    \reg_mstatus_prv_reg[1]_2 ,
    \bypass_mux_1_reg[36]_2 ,
    \bypass_mux_1_reg[38]_3 ,
    dcacheArb_io_requestor_1_req_bits_addr,
    \ex_ctrl_alu_fn_reg[3]_0 ,
    ex_reg_rvc_reg_2,
    ex_reg_rvc_reg_3,
    ex_reg_rvc_reg_4,
    \ex_ctrl_alu_fn_reg[3]_1 ,
    \ex_ctrl_alu_fn_reg[3]_2 ,
    \ex_ctrl_alu_fn_reg[3]_3 ,
    \ex_ctrl_alu_fn_reg[3]_4 ,
    \ex_reg_inst_reg[26]_0 ,
    ex_reg_rvc_reg_5,
    ex_reg_rvc_reg_6,
    ex_reg_rvc_reg_7,
    ex_reg_rvc_reg_8,
    ex_reg_rvc_reg_9,
    ex_reg_rvc_reg_10,
    ex_reg_rvc_reg_11,
    ex_reg_rvc_reg_12,
    ex_reg_rvc_reg_13,
    ex_reg_rvc_reg_14,
    ex_reg_rvc_reg_15,
    ex_reg_rvc_reg_16,
    ex_ctrl_alu_dw_reg_33,
    \ex_reg_inst_reg[10]_1 ,
    \ex_reg_inst_reg[10]_2 ,
    \ex_reg_inst_reg[10]_3 ,
    \ex_reg_inst_reg[10]_4 ,
    \ex_reg_inst_reg[10]_5 ,
    \ex_reg_inst_reg[10]_6 ,
    \ex_reg_inst_reg[10]_7 ,
    \ex_ctrl_alu_fn_reg[3]_5 ,
    \ex_ctrl_alu_fn_reg[3]_6 ,
    \ex_ctrl_alu_fn_reg[3]_7 ,
    \ex_ctrl_alu_fn_reg[3]_8 ,
    \ex_reg_pc_reg[39]_1 ,
    \ex_ctrl_alu_fn_reg[3]_9 );
  output req_dw_reg;
  output _T_1790;
  output mem_ctrl_mem;
  output mem_ctrl_fp;
  output wb_ctrl_mem;
  output ex_ctrl_jalr;
  output ex_reg_flush_pipe;
  output ex_ctrl_wxd;
  output ex_ctrl_div;
  output mem_reg_valid;
  output ex_reg_xcpt_interrupt;
  output mem_reg_xcpt_interrupt;
  output wb_ctrl_wxd;
  output mem_ctrl_jalr;
  output mem_ctrl_jal;
  output mem_reg_rvc;
  output mem_reg_rvc_reg_0;
  output ex_reg_xcpt;
  output mem_reg_xcpt;
  output wb_reg_xcpt;
  output wb_reg_replay;
  output wb_reg_valid;
  output wb_ctrl_div;
  output ex_reg_valid;
  output mem_ctrl_branch;
  output _T_1844;
  output mem_reg_sfence;
  output ex_ctrl_fence_i;
  output wb_ctrl_fence_i_reg_0;
  output mem_reg_flush_pipe;
  output \trig_pc_reg[0]_0 ;
  output mem_reg_slow_bypass;
  output ex_reg_rs_bypass_0_reg_0;
  output [34:0]_T_4899;
  output \reg_mtvec_reg[20] ;
  output \reg_mtvec_reg[21] ;
  output \reg_mtvec_reg[22] ;
  output reg_dcsr_step;
  output [5:0]_T_5044;
  output csr_io_bp_0_control_u;
  output csr_io_bp_0_control_s;
  output csr_io_bp_0_control_m;
  output csr_io_bp_0_control_action;
  output \_T_294_reg[3] ;
  output [0:0]\_T_281_reg[3] ;
  output csr_io_status_debug;
  output reg_mstatus_spie_reg;
  output reg_mstatus_mpie_reg;
  output dcache_io_ptw_status_sum;
  output dcache_io_ptw_status_mxr;
  output reg_singleStepped;
  output frontend_io_ptw_pmp_1_cfg_w;
  output [2:0]D;
  output buf__replay;
  output \ex_ctrl_sel_alu2_reg[1]_0 ;
  output buf__xcpt_ae_inst;
  output [0:0]_T_100;
  output \remainder_reg[129] ;
  output \remainder_reg[129]_0 ;
  output [0:0]_T_216;
  output \state_reg[2] ;
  output [0:0]Q;
  output \count_reg[0] ;
  output resHi_reg;
  output [64:0]\remainder_reg[65] ;
  output [66:0]\ex_reg_rs_msb_1_reg[29]_0 ;
  output \remainder_reg[31] ;
  output \remainder_reg[59] ;
  output [18:0]\s1_req_addr_reg[39] ;
  output [0:0]O;
  output [5:0]\divisor_reg[57] ;
  output \remainder_reg[33] ;
  output \remainder_reg[34] ;
  output \remainder_reg[35] ;
  output \remainder_reg[36] ;
  output \remainder_reg[37] ;
  output \remainder_reg[38] ;
  output \remainder_reg[39] ;
  output \remainder_reg[41] ;
  output \remainder_reg[42] ;
  output \remainder_reg[43] ;
  output \remainder_reg[44] ;
  output \remainder_reg[46] ;
  output \remainder_reg[47] ;
  output \remainder_reg[49] ;
  output \remainder_reg[50] ;
  output \remainder_reg[51] ;
  output \remainder_reg[52] ;
  output \remainder_reg[54] ;
  output \remainder_reg[55] ;
  output \remainder_reg[57] ;
  output \remainder_reg[58] ;
  output \remainder_reg[60] ;
  output \remainder_reg[61] ;
  output \remainder_reg[62] ;
  output neg_out_reg;
  output [19:0]\ex_reg_rs_msb_0_reg[27]_0 ;
  output \remainder_reg[63] ;
  output [3:0]\remainder_reg[107] ;
  output [3:0]\remainder_reg[111] ;
  output [3:0]\remainder_reg[115] ;
  output [3:0]\remainder_reg[119] ;
  output [0:0]\remainder_reg[127] ;
  output [3:0]\remainder_reg[127]_0 ;
  output [3:0]\remainder_reg[127]_1 ;
  output [3:0]\remainder_reg[127]_2 ;
  output [1:0]\remainder_reg[127]_3 ;
  output [3:0]\remainder_reg[123] ;
  output [3:0]\remainder_reg[127]_4 ;
  output [3:0]\remainder_reg[127]_5 ;
  output [2:0]\remainder_reg[129]_1 ;
  output [0:0]CO;
  output [3:0]\remainder_reg[91] ;
  output [3:0]\remainder_reg[95] ;
  output [3:0]\remainder_reg[99] ;
  output [3:0]\remainder_reg[103] ;
  output [0:0]\remainder_reg[115]_0 ;
  output [0:0]\remainder_reg[103]_0 ;
  output [2:0]\remainder_reg[103]_1 ;
  output [3:0]\remainder_reg[107]_0 ;
  output [3:0]\remainder_reg[111]_0 ;
  output [0:0]\remainder_reg[127]_6 ;
  output [2:0]\remainder_reg[115]_1 ;
  output [2:0]\reg_entries_0_reg[6] ;
  output [28:0]\reg_mtvec_reg[29] ;
  output \reg_entries_0_reg[0] ;
  output [2:0]\reg_entries_0_reg[6]_0 ;
  output [29:0]\reg_mtvec_reg[29]_0 ;
  output [1:0]\s2_req_addr_reg[31] ;
  output \reg_entries_0_reg[6]_1 ;
  output [27:0]\reg_mtvec_reg[29]_1 ;
  output [29:0]\reg_mtvec_reg[29]_2 ;
  output \reg_entries_0_reg[6]_2 ;
  output \reg_entries_0_reg[6]_3 ;
  output \reg_entries_0_reg[6]_4 ;
  output [29:0]\reg_mtvec_reg[29]_3 ;
  output \valid_reg[3] ;
  output frontend_io_cpu_sfence_valid;
  output [27:0]\reg_mtvec_reg[29]_4 ;
  output [28:0]\reg_mtvec_reg[29]_5 ;
  output [28:0]\reg_mtvec_reg[29]_6 ;
  output \reg_entries_1_reg[0] ;
  output \reg_entries_1_reg[0]_0 ;
  output \reg_entries_1_reg[0]_1 ;
  output \reg_entries_1_reg[0]_2 ;
  output \reg_entries_1_reg[0]_3 ;
  output \reg_entries_1_reg[0]_4 ;
  output \reg_entries_1_reg[0]_5 ;
  output \reg_entries_1_reg[0]_6 ;
  output s1_valid_reg;
  output mem_reg_replay_reg_0;
  output \reg_entries_1_reg[0]_7 ;
  output dcache_io_ptw_resp_bits_homogeneous;
  output [0:0]\reg_sbadaddr_reg[39] ;
  output [23:0]\reg_sscratch_reg[62] ;
  output [2:0]\reg_entries_1_reg[0]_8 ;
  output invalidated_reg;
  output [0:0]SR;
  output [0:0]\valid_reg[3]_0 ;
  output [0:0]\valid_reg[3]_1 ;
  output [0:0]\valid_reg[3]_2 ;
  output \valid_reg[3]_3 ;
  output \valid_reg[1] ;
  output \reg_entries_1_reg[0]_9 ;
  output [0:0]\reg_entries_0_reg[5] ;
  output _T_1081;
  output [1:0]frontend_io_ptw_status_prv;
  output [3:0]\reg_entries_0_reg[5]_0 ;
  output [0:0]\reg_pmp_5_cfg_a_reg[1] ;
  output [2:0]\reg_entries_1_reg[0]_10 ;
  output [3:0]\reg_entries_0_reg[5]_1 ;
  output [0:0]\reg_pmp_4_cfg_a_reg[1] ;
  output [2:0]\reg_entries_1_reg[0]_11 ;
  output [3:0]\reg_entries_0_reg[5]_2 ;
  output [3:0]\reg_entries_0_reg[5]_3 ;
  output [1:0]frontend_io_ptw_pmp_7_cfg_a;
  output [2:0]\reg_entries_1_reg[0]_12 ;
  output [3:0]\reg_entries_0_reg[5]_4 ;
  output [1:0]frontend_io_ptw_pmp_6_cfg_a;
  output [2:0]\reg_entries_1_reg[0]_13 ;
  output [3:0]\reg_entries_0_reg[5]_5 ;
  output [1:0]frontend_io_ptw_pmp_2_cfg_a;
  output [3:0]\reg_entries_0_reg[5]_6 ;
  output [1:0]frontend_io_ptw_pmp_1_cfg_a;
  output [2:0]\reg_entries_1_reg[0]_14 ;
  output [3:0]\reg_entries_0_reg[5]_7 ;
  output s2_valid_reg;
  output [0:0]frontend_io_ptw_ptbr_mode;
  output bad_va;
  output s2_tlb_resp_cacheable_reg;
  output [2:0]\reg_entries_0_reg[5]_8 ;
  output [2:0]\reg_entries_0_reg[5]_9 ;
  output [2:0]\reg_entries_0_reg[5]_10 ;
  output [2:0]\reg_entries_0_reg[5]_11 ;
  output [2:0]\reg_entries_0_reg[5]_12 ;
  output [2:0]\reg_entries_0_reg[5]_13 ;
  output [2:0]\reg_entries_0_reg[5]_14 ;
  output [2:0]\reg_entries_0_reg[5]_15 ;
  output [3:0]\reg_entries_0_reg[5]_16 ;
  output [3:0]\reg_entries_0_reg[5]_17 ;
  output [3:0]\reg_entries_0_reg[5]_18 ;
  output [3:0]\reg_entries_0_reg[5]_19 ;
  output [3:0]\reg_entries_0_reg[5]_20 ;
  output [3:0]\reg_entries_0_reg[5]_21 ;
  output [3:0]\reg_entries_0_reg[5]_22 ;
  output [3:0]\reg_entries_0_reg[5]_23 ;
  output [0:0]\reg_entries_0_reg[0]_0 ;
  output p_13_in;
  output [3:0]\reg_entries_0_reg[5]_24 ;
  output [3:0]\reg_entries_0_reg[5]_25 ;
  output [0:0]\reg_entries_0_reg[5]_26 ;
  output [3:0]\reg_entries_0_reg[5]_27 ;
  output [3:0]\reg_entries_0_reg[5]_28 ;
  output [0:0]\reg_entries_0_reg[5]_29 ;
  output [3:0]\reg_entries_0_reg[5]_30 ;
  output [3:0]\reg_entries_0_reg[5]_31 ;
  output [0:0]\reg_entries_0_reg[5]_32 ;
  output [3:0]\reg_entries_0_reg[5]_33 ;
  output [3:0]\reg_entries_0_reg[5]_34 ;
  output [0:0]\reg_entries_0_reg[5]_35 ;
  output [3:0]\reg_entries_0_reg[5]_36 ;
  output [3:0]\reg_entries_0_reg[5]_37 ;
  output [0:0]\reg_entries_0_reg[5]_38 ;
  output [3:0]\reg_entries_0_reg[5]_39 ;
  output [3:0]\reg_entries_0_reg[5]_40 ;
  output [0:0]\reg_entries_0_reg[5]_41 ;
  output [3:0]\reg_entries_0_reg[5]_42 ;
  output [3:0]\reg_entries_0_reg[5]_43 ;
  output [0:0]\reg_entries_0_reg[5]_44 ;
  output [3:0]\reg_entries_0_reg[5]_45 ;
  output [3:0]\reg_entries_0_reg[5]_46 ;
  output [0:0]\reg_entries_0_reg[5]_47 ;
  output [0:0]\reg_entries_0_reg[0]_1 ;
  output [0:0]\reg_entries_0_reg[0]_2 ;
  output [0:0]\reg_entries_0_reg[0]_3 ;
  output [0:0]\reg_entries_0_reg[0]_4 ;
  output [0:0]\reg_entries_0_reg[0]_5 ;
  output [0:0]\reg_entries_0_reg[0]_6 ;
  output [0:0]\reg_entries_0_reg[0]_7 ;
  output \ex_ctrl_sel_alu2_reg[1]_1 ;
  output \ex_ctrl_sel_alu2_reg[1]_2 ;
  output \ex_ctrl_sel_alu2_reg[1]_3 ;
  output _T_5074;
  output \_T_294_reg[0] ;
  output reg_mip_seip_reg;
  output \reg_pmp_7_addr_reg[29] ;
  output \reg_mtvec_reg[12] ;
  output [2:0]\reg_sscratch_reg[59] ;
  output \_T_1883_reg[1] ;
  output \reg_mbadaddr_reg[12] ;
  output [0:0]\reg_mie_reg[7] ;
  output \mem_reg_rs2_reg[7]_0 ;
  output [0:0]\s1_pc_reg[4] ;
  output \mem_reg_rs2_reg[6]_0 ;
  output \reg_sepc_reg[12] ;
  output \reg_mtvec_reg[8] ;
  output \reg_mepc_reg[12] ;
  output reg_mip_seip_reg_0;
  output [0:0]\s1_pc_reg[4]_0 ;
  output \reg_mtvec_reg[10] ;
  output \reg_mtvec_reg[11] ;
  output \reg_mtvec_reg[13] ;
  output [4:0]\reg_sscratch_reg[45] ;
  output [19:0]\r_pte_ppn_reg[19] ;
  output \reg_mtvec_reg[14] ;
  output \reg_mtvec_reg[15] ;
  output \reg_mtvec_reg[16] ;
  output \reg_mtvec_reg[17] ;
  output \reg_mtvec_reg[18] ;
  output \reg_mtvec_reg[19] ;
  output \reg_mtvec_reg[20]_0 ;
  output \reg_dpc_reg[12] ;
  output \reg_mtvec_reg[21]_0 ;
  output \reg_mtvec_reg[22]_0 ;
  output \reg_mtvec_reg[23] ;
  output \reg_mtvec_reg[24] ;
  output \reg_mtvec_reg[25] ;
  output \reg_mtvec_reg[26] ;
  output \reg_mtvec_reg[27] ;
  output \reg_mtvec_reg[28] ;
  output \reg_mtvec_reg[29]_7 ;
  output \reg_dscratch_reg[0] ;
  output \mem_reg_rs2_reg[0]_0 ;
  output \mem_reg_rs2_reg[1]_0 ;
  output [1:0]\reg_misa_reg[12] ;
  output \mem_reg_rs2_reg[2]_0 ;
  output \reg_mcause_reg[0] ;
  output \mem_reg_rs2_reg[3]_0 ;
  output \mem_reg_rs2_reg[4]_0 ;
  output \mem_reg_rs2_reg[5]_0 ;
  output [0:0]csr_io_tval;
  output \reg_stvec_reg[38] ;
  output \reg_stvec_reg[37] ;
  output \reg_stvec_reg[36] ;
  output \reg_stvec_reg[35] ;
  output \reg_stvec_reg[34] ;
  output \reg_stvec_reg[33] ;
  output \reg_stvec_reg[32] ;
  output \reg_mtvec_reg[31] ;
  output \reg_mtvec_reg[30] ;
  output \reg_sscratch_reg[0] ;
  output [13:0]\reg_bp_0_control_tmatch_reg[1] ;
  output \reg_sbadaddr_reg[0] ;
  output [0:0]\ex_cause_reg[1]_0 ;
  output \reg_misa_reg[0] ;
  output \reg_scause_reg[0] ;
  output \reg_pmp_2_addr_reg[29] ;
  output \_T_294_reg[0]_0 ;
  output reg_mstatus_mie;
  output reg_mstatus_mie_reg;
  output \reg_sscratch_reg[45]_0 ;
  output \reg_sptbr_ppn_reg[0] ;
  output \_T_1883_reg[0] ;
  output reg_debug_reg;
  output \reg_mstatus_prv_reg[1] ;
  output reg_mstatus_mpie_reg_0;
  output \reg_mstatus_mpp_reg[1] ;
  output \reg_mstatus_mpp_reg[0] ;
  output reg_mstatus_mie_reg_0;
  output \reg_dcsr_cause_reg[1] ;
  output \reg_scause_reg[1] ;
  output \s1_pc_reg[5] ;
  output \reg_scause_reg[3] ;
  output \reg_scause_reg[0]_0 ;
  output \reg_dcsr_cause_reg[0] ;
  output reg_wfi_reg;
  output \reg_scause_reg[1]_0 ;
  output reg_dcsr_prv;
  output \reg_bp_0_control_tmatch_reg[1]_0 ;
  output [0:0]\reg_scause_reg[2] ;
  output \reg_sepc_reg[26] ;
  output _T_481;
  output dcacheArb_io_requestor_1_req_valid;
  output [4:0]\s1_req_cmd_reg[4] ;
  output \state_reg[1] ;
  output [0:0]\s1_pc_reg[1] ;
  output [37:0]\s1_pc_reg[39]_0 ;
  output ibuf_io_inst_0_bits_xcpt0_ae_inst;
  output [19:0]\ex_reg_pc_reg[39]_0 ;
  output \ex_ctrl_sel_alu2_reg[1]_4 ;
  output ex_ctrl_mem_reg_0;
  output id_reg_fence_reg_0;
  output ex_ctrl_mem_reg_1;
  output ex_reg_rs_bypass_1_reg_0;
  output \ex_reg_rs_lsb_0_reg[0]_0 ;
  output \_T_2547_reg[1]_0 ;
  output ex_ctrl_mem_reg_2;
  output \ex_ctrl_sel_alu2_reg[1]_5 ;
  output ex_ctrl_mem_reg_3;
  output ex_ctrl_mem_reg_4;
  output ex_ctrl_mem_reg_5;
  output _T_1829;
  output \ex_reg_rs_lsb_0_reg[0]_1 ;
  output [24:0]\wb_reg_inst_reg[31]_0 ;
  output ex_ctrl_mem_reg_6;
  output \ex_reg_rs_lsb_0_reg[1]_0 ;
  output [62:0]_T_1406;
  output [43:0]_GEN_274;
  output [0:0]\_T_2547_reg[16]_0 ;
  output ex_ctrl_mem_reg_7;
  output ex_ctrl_mem_reg_8;
  output ex_ctrl_mem_reg_9;
  output [7:0]\mem_reg_inst_reg[31]_0 ;
  output \ex_reg_rs_msb_1_reg[61]_0 ;
  output [1:0]_T_1416;
  output p_31_in;
  output [2:0]\ex_reg_rs_msb_1_reg[61]_1 ;
  output ex_reg_rvc_reg_0;
  output _T_134;
  output \ex_reg_rs_msb_0_reg[10]_0 ;
  output \ex_reg_rs_msb_0_reg[8]_0 ;
  output \ex_reg_rs_msb_0_reg[9]_0 ;
  output \ex_reg_rs_msb_0_reg[11]_0 ;
  output \ex_reg_rs_msb_0_reg[12]_0 ;
  output \ex_reg_rs_msb_0_reg[13]_0 ;
  output \ex_reg_rs_msb_0_reg[14]_0 ;
  output \ex_reg_rs_msb_0_reg[15]_0 ;
  output \ex_reg_rs_msb_0_reg[16]_0 ;
  output \ex_reg_rs_msb_0_reg[17]_0 ;
  output \ex_reg_rs_msb_0_reg[18]_0 ;
  output \ex_reg_rs_msb_0_reg[19]_0 ;
  output \ex_reg_rs_msb_0_reg[20]_0 ;
  output \ex_reg_rs_msb_0_reg[21]_0 ;
  output \ex_reg_rs_msb_0_reg[22]_0 ;
  output \ex_reg_rs_msb_0_reg[23]_0 ;
  output \ex_reg_rs_msb_0_reg[24]_0 ;
  output \ex_reg_rs_msb_0_reg[25]_0 ;
  output \ex_reg_rs_msb_0_reg[26]_0 ;
  output \ex_reg_rs_msb_0_reg[27]_1 ;
  output [38:0]\reg_dpc_reg[39] ;
  output mem_reg_valid_reg_0;
  output dcacheArb_io_requestor_1_s1_kill;
  output frontend_io_cpu_req_bits_speculative;
  output \wb_reg_cause_reg[0]_0 ;
  output [1:0]\wb_reg_cause_reg[3]_0 ;
  output \ex_reg_rs_msb_1_reg[61]_2 ;
  output [4:0]\_T_2547_reg[31]_0 ;
  output \bypass_mux_2_reg[38]_0 ;
  output [1:0]\mem_reg_rs2_reg[3]_1 ;
  output [2:0]\reg_sbadaddr_reg[30] ;
  output [2:0]\reg_sbadaddr_reg[30]_0 ;
  output [2:0]\reg_sbadaddr_reg[30]_1 ;
  output [1:0]\reg_sbadaddr_reg[30]_2 ;
  output \lrscCount_reg[0] ;
  output \lrscCount_reg[0]_0 ;
  output \trig_state_reg[1]_0 ;
  output \trig_state_reg[0]_0 ;
  output \trig_state_reg[1]_1 ;
  output \trig_state_reg[1]_2 ;
  output \trig_pc_reg[0]_1 ;
  output trig_pc_valid_reg_0;
  output [3:0]\wb_reg_pc_reg[34]_0 ;
  output \bypass_mux_2_reg[35]_0 ;
  output [3:0]\bypass_mux_2_reg[31]_0 ;
  output ex_ctrl_mem_reg_10;
  output _T_1573;
  output ex_ctrl_mem_reg_11;
  output ex_sfence;
  output mem_reg_sfence_reg_0;
  output \trig_jalr_count_reg[0]_0 ;
  output [63:0]\a_data_reg[63] ;
  output [3:0]\s1_pc_reg[39]_1 ;
  output [3:0]\s1_pc_reg[39]_2 ;
  output [3:0]\s1_pc_reg[39]_3 ;
  output [3:0]\s1_pc_reg[39]_4 ;
  output [3:0]\trig_state_reg[1]_3 ;
  output [1:0]\trig_mem_data_reg[126]_0 ;
  output [3:0]\trig_state_reg[1]_4 ;
  output [3:0]\trig_state_reg[1]_5 ;
  output [3:0]\trig_state_reg[1]_6 ;
  output [3:0]\trig_state_reg[1]_7 ;
  output [0:0]\trig_state_reg[1]_8 ;
  output [3:0]\trig_jalr_count_reg[0]_1 ;
  output [3:0]\trig_jalr_count_reg[0]_2 ;
  output [3:0]\trig_jalr_count_reg[0]_3 ;
  output [3:0]\trig_jalr_count_reg[0]_4 ;
  output [3:0]\trig_jalr_count_reg[0]_5 ;
  output [0:0]\trig_jalr_count_reg[0]_6 ;
  output [3:0]\trig_pc_reg[0]_2 ;
  output [63:0]\trig_pc_reg[63]_0 ;
  output [32:0]\wb_reg_pc_reg[39]_0 ;
  output [3:0]\trig_pc_reg[0]_3 ;
  output [3:0]\trig_pc_reg[0]_4 ;
  output [3:0]\trig_pc_reg[0]_5 ;
  output [3:0]\trig_pc_reg[0]_6 ;
  output [0:0]\trig_pc_reg[0]_7 ;
  output [3:0]\s1_req_addr_reg[39]_0 ;
  output [3:0]\s1_req_addr_reg[39]_1 ;
  output [62:0]alu_io_in1;
  output [0:0]\mem_reg_pc_reg[31]_0 ;
  output \ex_ctrl_sel_alu1_reg[1]_0 ;
  output \ex_ctrl_sel_alu1_reg[0]_0 ;
  output \remainder_reg[33]_0 ;
  output \remainder_reg[34]_0 ;
  output \remainder_reg[35]_0 ;
  output \remainder_reg[36]_0 ;
  output \remainder_reg[37]_0 ;
  output \remainder_reg[38]_0 ;
  output [3:0]\s1_req_addr_reg[39]_2 ;
  output [3:0]\s1_req_addr_reg[39]_3 ;
  output [0:0]\reg_sbadaddr_reg[39]_0 ;
  output [3:0]\reg_sbadaddr_reg[39]_1 ;
  output [3:0]\reg_sbadaddr_reg[39]_2 ;
  output [0:0]\s1_pc_reg[39]_5 ;
  output mem_reg_slow_bypass_reg_0;
  output [2:0]dcacheArb_io_requestor_1_req_bits_typ;
  output [62:0]alu_io_in2;
  output [1:0]ex_ctrl_sel_alu2;
  output \mem_reg_rs2_reg[25]_0 ;
  output \bypass_mux_1_reg[6]_0 ;
  output \bypass_mux_1_reg[4]_0 ;
  output \reg_sbadaddr_reg[30]_3 ;
  output [2:0]\bypass_mux_1_reg[6]_1 ;
  output \bypass_mux_1_reg[0]_0 ;
  output [2:0]\reg_sbadaddr_reg[30]_4 ;
  output [0:0]\s1_req_addr_reg[3] ;
  output [0:0]\s1_req_addr_reg[39]_4 ;
  output [1:0]\reg_sbadaddr_reg[30]_5 ;
  output [2:0]\reg_sbadaddr_reg[30]_6 ;
  output [1:0]\reg_sbadaddr_reg[30]_7 ;
  output [1:0]\reg_sbadaddr_reg[30]_8 ;
  output [1:0]\reg_sbadaddr_reg[30]_9 ;
  output [0:0]\_T_389_reg[7] ;
  output \reg_entries_1_reg[0]_15 ;
  output \reg_entries_1_reg[0]_16 ;
  output \reg_entries_1_reg[0]_17 ;
  output \reg_entries_1_reg[0]_18 ;
  output \reg_entries_1_reg[0]_19 ;
  output \reg_entries_1_reg[0]_20 ;
  output \reg_entries_1_reg[0]_21 ;
  output \reg_entries_1_reg[0]_22 ;
  output \reg_entries_1_reg[0]_23 ;
  output \reg_entries_1_reg[0]_24 ;
  output \reg_entries_1_reg[0]_25 ;
  output \reg_entries_1_reg[0]_26 ;
  output \reg_entries_1_reg[0]_27 ;
  output \reg_entries_1_reg[0]_28 ;
  output \reg_entries_1_reg[0]_29 ;
  output \reg_entries_1_reg[0]_30 ;
  output \reg_entries_1_reg[0]_31 ;
  output [0:0]\reg_entries_1_reg[0]_32 ;
  output [0:0]\reg_entries_1_reg[0]_33 ;
  output [0:0]\reg_entries_1_reg[0]_34 ;
  output [0:0]\reg_entries_1_reg[0]_35 ;
  output [0:0]\reg_entries_1_reg[0]_36 ;
  output [0:0]\reg_entries_1_reg[0]_37 ;
  output [0:0]\reg_entries_1_reg[0]_38 ;
  output [0:0]\reg_entries_1_reg[0]_39 ;
  output [0:0]\reg_entries_1_reg[0]_40 ;
  output [0:0]\reg_entries_1_reg[0]_41 ;
  output [0:0]\reg_entries_1_reg[0]_42 ;
  output [0:0]\reg_entries_1_reg[0]_43 ;
  output [0:0]\reg_entries_1_reg[0]_44 ;
  output [0:0]\reg_entries_1_reg[0]_45 ;
  output [0:0]\reg_entries_1_reg[0]_46 ;
  output [0:0]\reg_entries_1_reg[0]_47 ;
  output [1:0]\reg_entries_0_reg[6]_5 ;
  output \reg_entries_0_reg[4] ;
  output \reg_entries_0_reg[6]_6 ;
  output _T_4068_ae_ld_reg;
  output _T_4068_pf_ld_reg;
  output \valid_reg[0] ;
  output \r_refill_waddr_reg[0] ;
  output \_T_973_reg[1] ;
  output \reg_entries_0_reg[6]_7 ;
  output \reg_entries_0_reg[4]_0 ;
  output [2:0]\reg_entries_0_reg[4]_1 ;
  output [2:0]\reg_entries_0_reg[4]_2 ;
  output [2:0]\reg_entries_0_reg[6]_8 ;
  output [2:0]\reg_entries_0_reg[6]_9 ;
  output [2:0]\reg_entries_0_reg[6]_10 ;
  output [2:0]\reg_entries_0_reg[6]_11 ;
  output [2:0]\reg_entries_0_reg[6]_12 ;
  output [2:0]\reg_entries_0_reg[6]_13 ;
  output [0:0]\reg_entries_0_reg[6]_14 ;
  output [1:0]\reg_entries_0_reg[6]_15 ;
  output [1:0]\reg_entries_0_reg[6]_16 ;
  output [1:0]\reg_entries_0_reg[6]_17 ;
  output [1:0]\reg_entries_0_reg[4]_3 ;
  output [1:0]\reg_entries_0_reg[4]_4 ;
  output [3:0]\reg_entries_0_reg[6]_18 ;
  output [3:0]\reg_entries_0_reg[6]_19 ;
  output [3:0]\reg_entries_0_reg[6]_20 ;
  output [3:0]\reg_entries_0_reg[6]_21 ;
  output [3:0]\reg_entries_0_reg[6]_22 ;
  output [3:0]\reg_entries_0_reg[6]_23 ;
  output [3:0]\reg_entries_0_reg[6]_24 ;
  output [3:0]\reg_entries_0_reg[6]_25 ;
  output [3:0]\reg_entries_0_reg[6]_26 ;
  output [3:0]\reg_entries_0_reg[4]_5 ;
  output [3:0]\reg_entries_0_reg[4]_6 ;
  output [3:0]\reg_entries_0_reg[4]_7 ;
  output \reg_entries_0_reg[4]_8 ;
  output [3:0]\reg_entries_0_reg[4]_9 ;
  output [2:0]\reg_entries_0_reg[6]_27 ;
  output [3:0]\reg_entries_0_reg[6]_28 ;
  output [3:0]\reg_entries_0_reg[6]_29 ;
  output [3:0]\reg_entries_0_reg[6]_30 ;
  output [3:0]\reg_entries_0_reg[6]_31 ;
  output [3:0]\reg_entries_0_reg[6]_32 ;
  output [3:0]\reg_entries_0_reg[6]_33 ;
  output [3:0]\reg_entries_0_reg[6]_34 ;
  output [3:0]\reg_entries_0_reg[6]_35 ;
  output [3:0]\reg_entries_0_reg[6]_36 ;
  output [3:0]\reg_entries_0_reg[4]_10 ;
  output [3:0]\reg_entries_0_reg[4]_11 ;
  output [3:0]\reg_entries_0_reg[4]_12 ;
  output [3:0]\reg_entries_0_reg[6]_37 ;
  output [2:0]\reg_entries_0_reg[6]_38 ;
  output [3:0]\reg_entries_0_reg[6]_39 ;
  output [2:0]\reg_entries_0_reg[4]_13 ;
  output [2:0]\reg_entries_0_reg[6]_40 ;
  output [2:0]\reg_entries_0_reg[6]_41 ;
  output \reg_entries_0_reg[4]_14 ;
  output \reg_entries_0_reg[4]_15 ;
  output \reg_entries_0_reg[4]_16 ;
  output \reg_entries_0_reg[6]_42 ;
  output [3:0]\reg_entries_0_reg[6]_43 ;
  output [3:0]\reg_entries_0_reg[6]_44 ;
  output \reg_entries_0_reg[6]_45 ;
  output [3:0]\reg_entries_0_reg[6]_46 ;
  output [3:0]\reg_entries_0_reg[6]_47 ;
  output \reg_entries_0_reg[6]_48 ;
  output [3:0]\reg_entries_0_reg[6]_49 ;
  output [3:0]\reg_entries_0_reg[6]_50 ;
  output \reg_entries_0_reg[4]_17 ;
  output [3:0]\reg_entries_0_reg[6]_51 ;
  output [3:0]\reg_entries_0_reg[6]_52 ;
  output \reg_entries_0_reg[6]_53 ;
  output [3:0]\reg_entries_0_reg[6]_54 ;
  output [3:0]\reg_entries_0_reg[6]_55 ;
  output \reg_entries_0_reg[4]_18 ;
  output [3:0]\reg_entries_0_reg[6]_56 ;
  output [3:0]\reg_entries_0_reg[6]_57 ;
  output \reg_entries_0_reg[4]_19 ;
  output [3:0]\reg_entries_0_reg[4]_20 ;
  output [3:0]\reg_entries_0_reg[4]_21 ;
  output \reg_entries_0_reg[4]_22 ;
  output [3:0]\reg_entries_0_reg[4]_23 ;
  output [3:0]\reg_entries_0_reg[4]_24 ;
  output \reg_entries_0_reg[4]_25 ;
  output _T_4068_pf_ld_reg_0;
  output _T_4068_pf_st_reg;
  output _T_4068_pf_ld_reg_1;
  output _T_4068_pf_ld_reg_2;
  output _T_4068_pf_st_reg_0;
  output _T_4068_pf_ld_reg_3;
  output _T_4068_pf_st_reg_1;
  output [15:0]\ex_reg_inst_reg[11]_0 ;
  output [0:0]\ex_cause_reg[1]_1 ;
  output [2:0]\ex_cause_reg[1]_2 ;
  output [2:0]\ex_cause_reg[1]_3 ;
  output [3:0]\ex_cause_reg[1]_4 ;
  output [3:0]\ex_cause_reg[1]_5 ;
  output [3:0]\ex_cause_reg[1]_6 ;
  output [3:0]\ex_cause_reg[1]_7 ;
  output [3:0]\ex_cause_reg[1]_8 ;
  output [3:0]\ex_cause_reg[1]_9 ;
  output [3:0]\ex_cause_reg[1]_10 ;
  output [3:0]\ex_cause_reg[1]_11 ;
  output [3:0]\ex_cause_reg[1]_12 ;
  output [2:0]\ex_cause_reg[1]_13 ;
  output [2:0]\ex_cause_reg[1]_14 ;
  output [3:0]\wb_reg_cause_reg[0]_1 ;
  output [3:0]\wb_reg_cause_reg[0]_2 ;
  output [3:0]\wb_reg_cause_reg[0]_3 ;
  output [0:0]\wb_reg_cause_reg[0]_4 ;
  output [3:0]\wb_reg_cause_reg[0]_5 ;
  output [3:0]\wb_reg_cause_reg[0]_6 ;
  output [3:0]\wb_reg_cause_reg[0]_7 ;
  output [3:0]\wb_reg_cause_reg[0]_8 ;
  output [3:0]\wb_reg_cause_reg[0]_9 ;
  output [3:0]\wb_reg_cause_reg[0]_10 ;
  output [3:0]\wb_reg_cause_reg[0]_11 ;
  output [3:0]\wb_reg_cause_reg[0]_12 ;
  output [2:0]\wb_reg_cause_reg[0]_13 ;
  output [2:0]\wb_reg_cause_reg[0]_14 ;
  output _T_217;
  output \bypass_mux_1_reg[32]_0 ;
  output \bypass_mux_1_reg[33]_0 ;
  output \bypass_mux_1_reg[34]_0 ;
  output \bypass_mux_1_reg[35]_0 ;
  output \bypass_mux_1_reg[36]_0 ;
  output \bypass_mux_1_reg[37]_0 ;
  output \bypass_mux_1_reg[38]_0 ;
  output \bypass_mux_1_reg[39]_0 ;
  output \bypass_mux_1_reg[40]_0 ;
  output \bypass_mux_1_reg[41]_0 ;
  output \bypass_mux_1_reg[42]_0 ;
  output \bypass_mux_1_reg[43]_0 ;
  output \bypass_mux_1_reg[44]_0 ;
  output \bypass_mux_1_reg[45]_0 ;
  output \bypass_mux_1_reg[46]_0 ;
  output \bypass_mux_1_reg[47]_0 ;
  output \bypass_mux_1_reg[60]_0 ;
  output \bypass_mux_1_reg[61]_0 ;
  output \bypass_mux_1_reg[62]_0 ;
  output \bypass_mux_1_reg[63]_0 ;
  output \bypass_mux_1_reg[48]_0 ;
  output \bypass_mux_1_reg[49]_0 ;
  output \bypass_mux_1_reg[50]_0 ;
  output \bypass_mux_1_reg[51]_0 ;
  output \bypass_mux_1_reg[52]_0 ;
  output \bypass_mux_1_reg[53]_0 ;
  output \bypass_mux_1_reg[54]_0 ;
  output \bypass_mux_1_reg[55]_0 ;
  output \bypass_mux_1_reg[56]_0 ;
  output \bypass_mux_1_reg[57]_0 ;
  output \bypass_mux_1_reg[58]_0 ;
  output \bypass_mux_1_reg[59]_0 ;
  output [3:0]\bypass_mux_1_reg[1]_0 ;
  output [0:0]shamt;
  output \bypass_mux_1_reg[62]_1 ;
  output \bypass_mux_1_reg[61]_1 ;
  output \bypass_mux_1_reg[60]_1 ;
  output \bypass_mux_1_reg[59]_1 ;
  output \bypass_mux_1_reg[58]_1 ;
  output \bypass_mux_1_reg[57]_1 ;
  output \bypass_mux_1_reg[56]_1 ;
  output \bypass_mux_1_reg[55]_1 ;
  output \bypass_mux_1_reg[54]_1 ;
  output \bypass_mux_1_reg[53]_1 ;
  output \bypass_mux_1_reg[52]_1 ;
  output \bypass_mux_1_reg[51]_1 ;
  output \bypass_mux_1_reg[50]_1 ;
  output \bypass_mux_1_reg[49]_1 ;
  output \bypass_mux_1_reg[48]_1 ;
  output \bypass_mux_1_reg[48]_2 ;
  output \bypass_mux_1_reg[47]_1 ;
  output \bypass_mux_1_reg[47]_2 ;
  output [0:0]_T_121;
  output \bypass_mux_1_reg[46]_1 ;
  output \bypass_mux_1_reg[46]_2 ;
  output \bypass_mux_1_reg[45]_1 ;
  output \bypass_mux_1_reg[45]_2 ;
  output \bypass_mux_1_reg[44]_1 ;
  output \bypass_mux_1_reg[44]_2 ;
  output \bypass_mux_1_reg[43]_1 ;
  output \bypass_mux_1_reg[43]_2 ;
  output \bypass_mux_1_reg[42]_1 ;
  output \bypass_mux_1_reg[42]_2 ;
  output \bypass_mux_1_reg[41]_1 ;
  output \bypass_mux_1_reg[41]_2 ;
  output \bypass_mux_1_reg[40]_1 ;
  output \bypass_mux_1_reg[40]_2 ;
  output \bypass_mux_1_reg[39]_1 ;
  output \bypass_mux_1_reg[39]_2 ;
  output \bypass_mux_1_reg[38]_1 ;
  output \bypass_mux_1_reg[38]_2 ;
  output \bypass_mux_1_reg[37]_1 ;
  output \bypass_mux_1_reg[37]_2 ;
  output \bypass_mux_1_reg[36]_1 ;
  output \bypass_mux_1_reg[35]_1 ;
  output \bypass_mux_1_reg[35]_2 ;
  output \bypass_mux_1_reg[34]_1 ;
  output \bypass_mux_1_reg[34]_2 ;
  output \bypass_mux_1_reg[33]_1 ;
  output \bypass_mux_1_reg[29]_0 ;
  output \bypass_mux_1_reg[33]_2 ;
  output \bypass_mux_1_reg[35]_3 ;
  output \bypass_mux_1_reg[29]_1 ;
  output \bypass_mux_1_reg[34]_3 ;
  output \bypass_mux_1_reg[34]_4 ;
  output \bypass_mux_1_reg[33]_3 ;
  output \bypass_mux_1_reg[33]_4 ;
  output \bypass_mux_1_reg[29]_2 ;
  output \bypass_mux_1_reg[29]_3 ;
  output \bypass_mux_1_reg[29]_4 ;
  output \bypass_mux_1_reg[23]_0 ;
  output \bypass_mux_1_reg[22]_0 ;
  output \bypass_mux_1_reg[21]_0 ;
  output \bypass_mux_1_reg[20]_0 ;
  output \bypass_mux_1_reg[19]_0 ;
  output \bypass_mux_1_reg[18]_0 ;
  output \bypass_mux_1_reg[17]_0 ;
  output \bypass_mux_1_reg[50]_2 ;
  output \bypass_mux_1_reg[51]_2 ;
  output \bypass_mux_1_reg[52]_2 ;
  output \bypass_mux_1_reg[53]_2 ;
  output \bypass_mux_1_reg[54]_2 ;
  output \bypass_mux_1_reg[55]_2 ;
  output \bypass_mux_1_reg[56]_2 ;
  output \bypass_mux_1_reg[57]_2 ;
  output \bypass_mux_1_reg[58]_2 ;
  output \bypass_mux_1_reg[59]_2 ;
  output \bypass_mux_1_reg[3]_0 ;
  output \bypass_mux_1_reg[2]_0 ;
  output \bypass_mux_1_reg[1]_1 ;
  output \bypass_mux_1_reg[1]_2 ;
  output [0:0]mem_br_taken__reg_0;
  output \bypass_mux_1_reg[48]_3 ;
  output \bypass_mux_1_reg[49]_2 ;
  output \bypass_mux_1_reg[50]_3 ;
  output \bypass_mux_1_reg[51]_3 ;
  output \bypass_mux_1_reg[52]_3 ;
  output \bypass_mux_1_reg[53]_3 ;
  output \bypass_mux_1_reg[54]_3 ;
  output \bypass_mux_1_reg[55]_3 ;
  output \bypass_mux_1_reg[56]_3 ;
  output \bypass_mux_1_reg[57]_3 ;
  output \bypass_mux_1_reg[58]_3 ;
  output \bypass_mux_1_reg[59]_3 ;
  input host_clk;
  input id_ctrl_mem;
  input \buf__data_reg[1] ;
  input _T_1821;
  input id_ctrl_wxd;
  input \buf__data_reg[1]_0 ;
  input id_ctrl_jal;
  input mem_reg_xcpt0;
  input \buf__data_reg[1]_1 ;
  input id_ctrl_rxs2;
  input id_ctrl_fence_i;
  input ex_ctrl_div_reg_0;
  input mem_reg_flush_pipe_reg_0;
  input mem_reg_sfence_reg_1;
  input ex_reg_rvc_reg_1;
  input target_reset;
  input trig_pc_valid_reg_1;
  input mem_ctrl_fence_i_reg_0;
  input ex_ctrl_alu_dw_reg_0;
  input mem_reg_slow_bypass_reg_1;
  input ex_reg_rs_bypass_0_reg_1;
  input reg_debug_reg_0;
  input tile_auto_int_sync_xing_sinklzy_in_2_sync_0;
  input sys_reset_reg;
  input reg_debug_reg_1;
  input \ex_ctrl_csr_reg[2]_0 ;
  input \ex_ctrl_csr_reg[1]_0 ;
  input \ex_ctrl_csr_reg[0]_0 ;
  input buf__pc;
  input frontend_io_cpu_resp_bits_replay;
  input frontend_io_cpu_resp_bits_xcpt_pf_inst;
  input frontend_io_cpu_resp_bits_xcpt_ae_inst;
  input nBufValid_reg;
  input \state_reg[1]_0 ;
  input doUncachedResp_reg;
  input [0:0]\bypass_mux_2_reg[9]_0 ;
  input \state_reg[0] ;
  input [3:0]S;
  input [3:0]\remainder_reg[71] ;
  input [3:0]\remainder_reg[75] ;
  input [3:0]\remainder_reg[79] ;
  input [3:0]\remainder_reg[83] ;
  input [3:0]\remainder_reg[87] ;
  input [3:0]\remainder_reg[91]_0 ;
  input [3:0]\remainder_reg[95]_0 ;
  input [3:0]\remainder_reg[99]_0 ;
  input [3:0]\remainder_reg[103]_2 ;
  input [3:0]\remainder_reg[107]_1 ;
  input [3:0]\remainder_reg[111]_1 ;
  input [3:0]\remainder_reg[115]_2 ;
  input [3:0]\remainder_reg[119]_0 ;
  input [3:0]\remainder_reg[123]_0 ;
  input [3:0]\remainder_reg[127]_7 ;
  input [0:0]\remainder_reg[128] ;
  input [0:0]\divisor_reg[35] ;
  input [0:0]\divisor_reg[52] ;
  input [2:0]\remainder_reg[64] ;
  input [3:0]\remainder_reg[64]_0 ;
  input [3:0]\remainder_reg[64]_1 ;
  input [2:0]\remainder_reg[64]_2 ;
  input [0:0]\divisor_reg[1] ;
  input [0:0]\divisor_reg[18] ;
  input [2:0]\divisor_reg[15] ;
  input [3:0]\divisor_reg[15]_0 ;
  input [3:0]\divisor_reg[15]_1 ;
  input [3:0]\divisor_reg[15]_2 ;
  input [1:0]DI;
  input [3:0]\divisor_reg[15]_3 ;
  input [3:0]\divisor_reg[15]_4 ;
  input [3:0]\divisor_reg[15]_5 ;
  input [3:0]\divisor_reg[15]_6 ;
  input [3:0]\divisor_reg[15]_7 ;
  input [1:0]\divisor_reg[15]_8 ;
  input [2:0]\divisor_reg[32] ;
  input [2:0]\remainder_reg[64]_3 ;
  input [3:0]\remainder_reg[64]_4 ;
  input [3:0]\remainder_reg[64]_5 ;
  input [3:0]\remainder_reg[64]_6 ;
  input [3:0]\divisor_reg[51] ;
  input [3:0]\divisor_reg[32]_0 ;
  input [3:0]\divisor_reg[32]_1 ;
  input [0:0]\remainder_reg[64]_7 ;
  input [3:0]\remainder_reg[64]_8 ;
  input [0:0]\remainder_reg[64]_9 ;
  input [9:0]\reg_entries_4_reg[61] ;
  input [10:0]\s1_req_addr_reg[31] ;
  input dcache_io_ptw_resp_valid;
  input [19:0]\r_pte_ppn_reg[19]_0 ;
  input s1_req_phys_reg;
  input \reg_pmp_7_cfg_a_reg[0] ;
  input s2_replay;
  input \r_pte_ppn_reg[7] ;
  input \r_pte_ppn_reg[7]_0 ;
  input \r_pte_ppn_reg[7]_1 ;
  input \r_pte_ppn_reg[7]_2 ;
  input \r_pte_ppn_reg[7]_3 ;
  input \r_pte_ppn_reg[7]_4 ;
  input \r_pte_ppn_reg[7]_5 ;
  input \r_pte_ppn_reg[7]_6 ;
  input [0:0]io_mask;
  input dcache_io_ptw_resp_bits_ae;
  input \s1_req_typ_reg[1] ;
  input \r_pte_ppn_reg[5] ;
  input [12:0]_T_200__0;
  input [11:0]\s1_pc_reg[39]_6 ;
  input dcacheArb_io_requestor_1_s2_nack;
  input invalidated;
  input refill_valid;
  input p_2_in;
  input [0:0]_T_1432;
  input [0:0]\valid_reg[3]_4 ;
  input [0:0]\reg_entries_3_reg[11] ;
  input [1:0]\r_refill_waddr_reg[1] ;
  input \s1_pc_reg[31] ;
  input resp_valid_1_reg;
  input [0:0]\reg_pmp_0_addr_reg[28] ;
  input [0:0]_T_726;
  input [0:0]\reg_pmp_5_addr_reg[28] ;
  input [0:0]\reg_pmp_4_addr_reg[28] ;
  input [0:0]\reg_pmp_3_addr_reg[28] ;
  input [0:0]\reg_pmp_2_addr_reg[28] ;
  input [0:0]\reg_pmp_7_addr_reg[28] ;
  input [0:0]\reg_pmp_6_addr_reg[28] ;
  input [0:0]\reg_pmp_1_addr_reg[28] ;
  input hitsVec_4;
  input [0:0]_T_382;
  input \reg_pmp_0_addr_reg[29] ;
  input \reg_pmp_1_addr_reg[29] ;
  input \reg_pmp_2_addr_reg[29]_0 ;
  input \reg_pmp_6_addr_reg[29] ;
  input \reg_pmp_7_addr_reg[29]_0 ;
  input \reg_pmp_3_addr_reg[29] ;
  input \reg_pmp_4_addr_reg[29] ;
  input \reg_pmp_5_addr_reg[29] ;
  input [2:0]_T_382__0;
  input \s1_pc_reg[26] ;
  input \reg_pmp_5_addr_reg[17] ;
  input \reg_pmp_4_addr_reg[17] ;
  input \reg_pmp_3_addr_reg[17] ;
  input \reg_pmp_7_addr_reg[17] ;
  input \reg_pmp_6_addr_reg[17] ;
  input \reg_pmp_2_addr_reg[17] ;
  input \reg_pmp_1_addr_reg[17] ;
  input \reg_pmp_0_addr_reg[17] ;
  input [0:0]_T_480;
  input \reg_pmp_5_addr_reg[19] ;
  input \reg_pmp_4_addr_reg[19] ;
  input \reg_pmp_3_addr_reg[19] ;
  input \reg_pmp_7_addr_reg[19] ;
  input \reg_pmp_6_addr_reg[19] ;
  input \reg_pmp_2_addr_reg[19] ;
  input \reg_pmp_1_addr_reg[19] ;
  input \reg_pmp_0_addr_reg[19] ;
  input \reg_pmp_5_addr_reg[13] ;
  input \reg_pmp_4_addr_reg[13] ;
  input \reg_pmp_3_addr_reg[13] ;
  input \reg_pmp_7_addr_reg[13] ;
  input \reg_pmp_6_addr_reg[13] ;
  input \reg_pmp_2_addr_reg[13] ;
  input \reg_pmp_1_addr_reg[13] ;
  input \reg_pmp_0_addr_reg[13] ;
  input nBufValid_reg_0;
  input nBufValid_reg_1;
  input [1:0]frontend_io_cpu_resp_bits_data;
  input [0:0]ibuf_io_inst_0_bits_raw;
  input \wb_reg_inst_reg[21]_0 ;
  input \wb_reg_cause_reg[63]_0 ;
  input \wb_reg_inst_reg[21]_1 ;
  input \wb_reg_inst_reg[22]_0 ;
  input \wb_reg_inst_reg[21]_2 ;
  input \wb_reg_inst_reg[21]_3 ;
  input wb_reg_replay_reg_0;
  input \wb_ctrl_csr_reg[2]_0 ;
  input \wb_reg_inst_reg[29]_0 ;
  input tile_auto_int_sync_xing_sinklzy_in_0_sync_0;
  input \wb_reg_inst_reg[21]_4 ;
  input \wb_reg_inst_reg[21]_5 ;
  input \reg_pmp_5_addr_reg[20] ;
  input \wb_reg_inst_reg[30]_0 ;
  input \wb_reg_inst_reg[30]_1 ;
  input \reg_mstatus_prv_reg[1]_0 ;
  input tile_auto_int_sync_xing_sinklzy_in_0_sync_1;
  input tile_auto_int_sync_xing_sinklzy_in_1_sync_0;
  input \wb_reg_inst_reg[29]_1 ;
  input reg_debug_reg_2;
  input \wb_reg_inst_reg[22]_1 ;
  input \wb_reg_cause_reg[2]_0 ;
  input \wb_ctrl_csr_reg[0]_0 ;
  input dcache_io_cpu_invalidate_lr;
  input \wb_reg_inst_reg[26]_0 ;
  input \reg_mstatus_prv_reg[1]_1 ;
  input wb_reg_replay_reg_1;
  input [0:0]\_T_294_reg[0]_1 ;
  input [0:0]\_T_281_reg[0] ;
  input [0:0]q_reg;
  input \state_reg[0]_0 ;
  input \state_reg[1]_1 ;
  input \state_reg[0]_1 ;
  input [0:0]\s2_pc_reg[1] ;
  input [38:0]frontend_io_cpu_resp_bits_pc;
  input [18:0]\elts_0_pc_reg[39] ;
  input nBufValid_reg_2;
  input frontend_io_cpu_resp_valid;
  input buf__xcpt_pf_inst_reg;
  input reg_mstatus_tvm_reg;
  input \s2_req_tag_reg[5] ;
  input \wb_reg_inst_reg[7]_0 ;
  input \buf__data_reg[3] ;
  input dcacheArb_io_requestor_1_ordered;
  input \buf__data_reg[2] ;
  input nBufValid_reg_3;
  input \buf__data_reg[4] ;
  input nBufValid_reg_4;
  input [4:0]ibuf_io_inst_0_bits_inst_rs2;
  input \buf__data_reg[3]_0 ;
  input [4:0]ibuf_io_inst_0_bits_inst_rs1;
  input \_T_2547_reg[16]_1 ;
  input nBufValid_reg_5;
  input \ex_reg_inst_reg[10]_0 ;
  input \wb_reg_inst_reg[7]_1 ;
  input \state_reg[0]_2 ;
  input \buf__data_reg[12] ;
  input [1:0]_T_1005;
  input \mem_reg_inst_reg[11]_0 ;
  input [4:0]ibuf_io_inst_0_bits_inst_rd;
  input [19:0]\s2_req_typ_reg[0] ;
  input \req_tag_reg[4] ;
  input ex_ctrl_wxd_reg_0;
  input reg_bp_0_control_action_reg;
  input buf__xcpt_pf_inst_reg_0;
  input \s2_req_cmd_reg[1] ;
  input [43:0]dcacheArb_io_requestor_1_resp_bits_data;
  input \reg_mtvec_reg[4] ;
  input wb_reg_valid_reg_0;
  input dcacheArb_io_requestor_1_replay_next;
  input mem_reg_sfence_reg_2;
  input dcacheArb_io_requestor_1_resp_valid;
  input dcacheArb_io_requestor_1_req_ready;
  input wb_reg_replay_reg_2;
  input \s2_req_tag_reg[5]_0 ;
  input [4:0]\s2_req_tag_reg[6] ;
  input dcacheArb_io_requestor_1_resp_bits_replay;
  input \req_tag_reg[0] ;
  input \s2_req_tag_reg[6]_0 ;
  input \wb_reg_inst_reg[9]_0 ;
  input \req_tag_reg[1] ;
  input \wb_reg_inst_reg[9]_1 ;
  input \req_tag_reg[1]_0 ;
  input \wb_reg_inst_reg[9]_2 ;
  input \req_tag_reg[1]_1 ;
  input \req_tag_reg[0]_0 ;
  input \req_tag_reg[1]_2 ;
  input \req_tag_reg[1]_3 ;
  input \req_tag_reg[1]_4 ;
  input \wb_reg_inst_reg[9]_3 ;
  input [39:0]p_0_in;
  input dcacheArb_io_requestor_1_s2_xcpt_ma_st;
  input wb_ctrl_mem_reg_0;
  input dcacheArb_io_requestor_1_s2_xcpt_pf_st;
  input dcacheArb_io_requestor_1_s2_xcpt_pf_ld;
  input dcacheArb_io_requestor_1_s2_xcpt_ma_ld;
  input [0:0]\bypass_mux_2_reg[63]_0 ;
  input [0:0]\bypass_mux_2_reg[63]_1 ;
  input [0:0]\trig_mem_data_reg[127]_0 ;
  input [0:0]\trig_mem_data_reg[63]_0 ;
  input trig_pc_valid_reg_2;
  input [0:0]\bypass_mux_1_reg[63]_1 ;
  input [0:0]\bypass_mux_1_reg[63]_2 ;
  input \trig_state_reg[0]_1 ;
  input [0:0]\trig_pc_reg[63]_1 ;
  input [63:0]dcacheArb_io_requestor_1_resp_bits_data_word_bypass;
  input [1:0]\ex_ctrl_mem_type_reg[0]_0 ;
  input \ex_ctrl_sel_imm_reg[1]_0 ;
  input [0:0]\wb_reg_cause_reg[63]_1 ;
  input [0:0]\wb_reg_cause_reg[63]_2 ;
  input [0:0]\wb_reg_cause_reg[63]_3 ;
  input [0:0]\wb_reg_cause_reg[63]_4 ;
  input [0:0]\wb_reg_cause_reg[63]_5 ;
  input [0:0]\wb_reg_cause_reg[63]_6 ;
  input \ex_ctrl_sel_imm_reg[1]_1 ;
  input \reg_pmp_5_cfg_a_reg[1]_0 ;
  input \count_reg[1] ;
  input \r_pte_ppn_reg[3] ;
  input \r_pte_ppn_reg[5]_0 ;
  input \r_pte_ppn_reg[16] ;
  input \count_reg[1]_0 ;
  input \r_pte_ppn_reg[3]_0 ;
  input \r_pte_ppn_reg[5]_1 ;
  input \r_pte_ppn_reg[16]_0 ;
  input \r_pte_ppn_reg[3]_1 ;
  input \r_pte_ppn_reg[5]_2 ;
  input \r_pte_ppn_reg[16]_1 ;
  input \r_pte_ppn_reg[3]_2 ;
  input \r_pte_ppn_reg[5]_3 ;
  input \r_pte_ppn_reg[16]_2 ;
  input _T_1156;
  input \r_pte_ppn_reg[3]_3 ;
  input \r_pte_ppn_reg[5]_4 ;
  input \r_pte_ppn_reg[16]_3 ;
  input _T_931;
  input [0:0]\reg_pmp_0_addr_reg[28]_0 ;
  input \r_pte_ppn_reg[3]_4 ;
  input \r_pte_ppn_reg[5]_5 ;
  input \r_pte_ppn_reg[16]_4 ;
  input \count_reg[1]_1 ;
  input \r_pte_ppn_reg[3]_5 ;
  input \r_pte_ppn_reg[5]_6 ;
  input \r_pte_ppn_reg[16]_5 ;
  input \count_reg[1]_2 ;
  input \r_pte_ppn_reg[3]_6 ;
  input \r_pte_ppn_reg[5]_7 ;
  input \r_pte_ppn_reg[16]_6 ;
  input [1:0]dcache_io_ptw_resp_bits_level;
  input [0:0]\reg_pmp_5_addr_reg[28]_0 ;
  input [0:0]\reg_pmp_6_addr_reg[28]_0 ;
  input [0:0]\reg_pmp_1_addr_reg[28]_0 ;
  input [0:0]\reg_pmp_2_addr_reg[28]_0 ;
  input [0:0]\reg_pmp_7_addr_reg[28]_0 ;
  input [0:0]\reg_pmp_4_addr_reg[28]_0 ;
  input [0:0]\reg_pmp_3_addr_reg[28]_0 ;
  input s1_req_phys_reg_0;
  input \reg_entries_4_reg[61]_0 ;
  input \valid_reg[4] ;
  input [0:0]\reg_entries_0_reg[10] ;
  input \valid_reg[2] ;
  input \valid_reg[0]_0 ;
  input \valid_reg[1]_0 ;
  input \reg_pmp_1_cfg_a_reg[0] ;
  input \reg_pmp_2_cfg_a_reg[0] ;
  input resp_valid_0_reg;
  input reg_pmp_1_cfg_w_reg;
  input \s1_req_addr_reg[2] ;
  input \s1_req_typ_reg[0] ;
  input \s1_req_typ_reg[0]_0 ;
  input tlb_io_req_bits_sfence_bits_rs2;
  input [0:0]\reg_pmp_1_addr_reg[29]_0 ;
  input \s1_req_addr_reg[2]_0 ;
  input \r_pte_ppn_reg[11] ;
  input [0:0]_T_382_0;
  input \r_pte_ppn_reg[16]_7 ;
  input [0:0]\reg_pmp_3_addr_reg[29]_0 ;
  input \reg_pmp_2_addr_reg[0] ;
  input [0:0]\reg_pmp_2_addr_reg[29]_1 ;
  input \s1_req_typ_reg[0]_1 ;
  input \s1_req_typ_reg[0]_2 ;
  input \reg_pmp_4_addr_reg[14] ;
  input \reg_pmp_4_addr_reg[0] ;
  input [0:0]\reg_pmp_5_addr_reg[29]_0 ;
  input \s1_req_addr_reg[2]_1 ;
  input \s1_req_typ_reg[0]_3 ;
  input [0:0]\reg_pmp_4_addr_reg[29]_0 ;
  input \reg_pmp_3_addr_reg[23] ;
  input \reg_pmp_3_addr_reg[29]_1 ;
  input \r_pte_ppn_reg[15] ;
  input [0:0]\reg_pmp_6_addr_reg[29]_0 ;
  input \s1_req_addr_reg[2]_2 ;
  input [0:0]\reg_pmp_0_addr_reg[29]_0 ;
  input \reg_pmp_0_addr_reg[23] ;
  input \r_pte_ppn_reg[6] ;
  input [0:0]\reg_pmp_7_addr_reg[29]_1 ;
  input \r_pte_ppn_reg[10] ;
  input \r_pte_ppn_reg[3]_7 ;
  input \reg_pmp_7_addr_reg[23] ;
  input \reg_pmp_7_addr_reg[29]_2 ;
  input \r_pte_ppn_reg[2] ;
  input \r_pte_ppn_reg[14] ;
  input \r_pte_ppn_reg[7]_7 ;
  input \r_pte_ppn_reg[13] ;
  input \r_pte_ppn_reg[0] ;
  input \r_pte_ppn_reg[8] ;
  input \r_pte_ppn_reg[4] ;
  input \r_pte_ppn_reg[1] ;
  input \r_pte_ppn_reg[17] ;
  input \r_pte_ppn_reg[18] ;
  input [5:0]_T_1701;
  input \reg_pmp_7_addr_reg[17]_0 ;
  input \r_pte_ppn_reg[9] ;
  input \reg_pmp_3_addr_reg[18] ;
  input \r_pte_ppn_reg[12] ;
  input [2:0]\reg_entries_2_reg[12] ;
  input [0:0]\reg_entries_1_reg[12] ;
  input [2:0]\reg_entries_3_reg[12] ;
  input [24:0]\remainder_reg[62]_0 ;
  input sys_reset_reg_0;
  input [4:0]ADDRA;
  input [4:0]nBufValid_reg_6;
  input [4:0]_T_909;
  input [2:0]_T_1142;
  input [0:0]_T_877;
  input [14:0]_T_889;
  input [0:0]_T_1031;
  input [3:0]\buf__data_reg[3]_1 ;
  input ex_ctrl_alu_dw_reg_1;
  input ex_ctrl_alu_dw_reg_2;
  input ex_ctrl_alu_dw_reg_3;
  input ex_ctrl_alu_dw_reg_4;
  input ex_ctrl_alu_dw_reg_5;
  input ex_ctrl_alu_dw_reg_6;
  input ex_ctrl_alu_dw_reg_7;
  input ex_ctrl_alu_dw_reg_8;
  input ex_ctrl_alu_dw_reg_9;
  input ex_ctrl_alu_dw_reg_10;
  input ex_ctrl_alu_dw_reg_11;
  input ex_ctrl_alu_dw_reg_12;
  input ex_ctrl_alu_dw_reg_13;
  input ex_ctrl_alu_dw_reg_14;
  input ex_ctrl_alu_dw_reg_15;
  input ex_ctrl_alu_dw_reg_16;
  input ex_ctrl_alu_dw_reg_17;
  input ex_ctrl_alu_dw_reg_18;
  input ex_ctrl_alu_dw_reg_19;
  input ex_ctrl_alu_dw_reg_20;
  input ex_ctrl_alu_dw_reg_21;
  input ex_ctrl_alu_dw_reg_22;
  input ex_ctrl_alu_dw_reg_23;
  input ex_ctrl_alu_dw_reg_24;
  input ex_ctrl_alu_dw_reg_25;
  input ex_ctrl_alu_dw_reg_26;
  input ex_ctrl_alu_dw_reg_27;
  input ex_ctrl_alu_dw_reg_28;
  input ex_ctrl_alu_dw_reg_29;
  input ex_ctrl_alu_dw_reg_30;
  input ex_ctrl_alu_dw_reg_31;
  input ex_ctrl_alu_dw_reg_32;
  input \buf__data_reg[1]_2 ;
  input [0:0]E;
  input [1:0]\buf__data_reg[3]_2 ;
  input nBufValid_reg_7;
  input [1:0]ex_ctrl_wxd_reg_1;
  input [0:0]\mem_reg_inst_reg[9]_0 ;
  input [63:0]out;
  input mem_ctrl_branch_reg_0;
  input [1:0]\buf__data_reg[1]_3 ;
  input [0:0]\mem_reg_inst_reg[9]_1 ;
  input [61:0]\bypass_mux_2_reg[63]_2 ;
  input [3:0]\buf__data_reg[3]_3 ;
  input [1:0]mem_reg_xcpt_interrupt_reg_0;
  input [2:0]nBufValid_reg_8;
  input buf__xcpt_pf_inst_reg_1;
  input \buf__data_reg[4]_0 ;
  input elts_0_xcpt_ae_inst_reg;
  input buf__xcpt_pf_inst_reg_2;
  input \reg_misa_reg[12]_0 ;
  input [1:0]id_ctrl_sel_alu1;
  input sys_reset_reg_1;
  input sys_reset_reg_2;
  input [0:0]\wb_ctrl_csr_reg[0]_1 ;
  input [38:0]\wb_reg_pc_reg[39]_1 ;
  input [0:0]\wb_ctrl_csr_reg[0]_2 ;
  input [39:0]\wb_ctrl_csr_reg[0]_3 ;
  input [0:0]\wb_ctrl_csr_reg[0]_4 ;
  input [4:0]\wb_ctrl_csr_reg[0]_5 ;
  input [0:0]\wb_ctrl_csr_reg[0]_6 ;
  input [38:0]\wb_reg_pc_reg[39]_2 ;
  input [0:0]\wb_ctrl_csr_reg[0]_7 ;
  input [5:0]\wb_ctrl_csr_reg[0]_8 ;
  input [0:0]\wb_ctrl_csr_reg[0]_9 ;
  input [38:0]\wb_reg_pc_reg[39]_3 ;
  input \wb_ctrl_csr_reg[0]_10 ;
  input [0:0]nBufValid_reg_9;
  input [15:0]\elts_0_data_reg[15] ;
  input \reg_bp_0_address_reg[3] ;
  input [0:0]\reg_bp_0_address_reg[36] ;
  input [0:0]\elts_0_pc_reg[38] ;
  input \reg_mstatus_prv_reg[1]_2 ;
  input [0:0]\bypass_mux_1_reg[36]_2 ;
  input [0:0]\bypass_mux_1_reg[38]_3 ;
  input [32:0]dcacheArb_io_requestor_1_req_bits_addr;
  input \ex_ctrl_alu_fn_reg[3]_0 ;
  input ex_reg_rvc_reg_2;
  input ex_reg_rvc_reg_3;
  input ex_reg_rvc_reg_4;
  input \ex_ctrl_alu_fn_reg[3]_1 ;
  input \ex_ctrl_alu_fn_reg[3]_2 ;
  input \ex_ctrl_alu_fn_reg[3]_3 ;
  input \ex_ctrl_alu_fn_reg[3]_4 ;
  input \ex_reg_inst_reg[26]_0 ;
  input ex_reg_rvc_reg_5;
  input ex_reg_rvc_reg_6;
  input ex_reg_rvc_reg_7;
  input ex_reg_rvc_reg_8;
  input ex_reg_rvc_reg_9;
  input ex_reg_rvc_reg_10;
  input ex_reg_rvc_reg_11;
  input ex_reg_rvc_reg_12;
  input ex_reg_rvc_reg_13;
  input ex_reg_rvc_reg_14;
  input ex_reg_rvc_reg_15;
  input ex_reg_rvc_reg_16;
  input ex_ctrl_alu_dw_reg_33;
  input \ex_reg_inst_reg[10]_1 ;
  input \ex_reg_inst_reg[10]_2 ;
  input \ex_reg_inst_reg[10]_3 ;
  input \ex_reg_inst_reg[10]_4 ;
  input \ex_reg_inst_reg[10]_5 ;
  input \ex_reg_inst_reg[10]_6 ;
  input \ex_reg_inst_reg[10]_7 ;
  input \ex_ctrl_alu_fn_reg[3]_5 ;
  input \ex_ctrl_alu_fn_reg[3]_6 ;
  input \ex_ctrl_alu_fn_reg[3]_7 ;
  input \ex_ctrl_alu_fn_reg[3]_8 ;
  input [0:0]\ex_reg_pc_reg[39]_1 ;
  input [0:0]\ex_ctrl_alu_fn_reg[3]_9 ;
  output [24:0]_T_2177;

  wire \<const0> ;
  wire \<const1> ;
  wire [4:0]ADDRA;
  wire [0:0]CO;
  wire [2:0]D;
  wire [1:0]DI;
  wire [0:0]E;
  wire [0:0]O;
  wire [0:0]Q;
  wire [3:0]S;
  wire [0:0]SR;
  wire [43:0]_GEN_274;
  wire [125:0]_GEN_277;
  wire [0:0]_T_100;
  wire [1:0]_T_1005;
  wire [0:0]_T_1031;
  wire _T_1081;
  wire [2:0]_T_1142;
  wire _T_1156;
  wire [0:0]_T_121;
  wire _T_134;
  wire [4:3]_T_1396__T_2475_addr;
  wire _T_1396_reg_r1_0_31_0_5_i_44_n_0;
  wire [62:0]_T_1406;
  wire [1:1]_T_1406_1;
  wire [1:0]_T_1416;
  wire [63:2]_T_1416_0;
  wire [0:0]_T_1432;
  wire _T_1573;
  wire [5:0]_T_1701;
  wire _T_1710;
  wire _T_1790;
  wire _T_1821;
  wire _T_1829;
  wire _T_1844;
  wire [61:0]_T_1856;
  wire _T_1865;
  wire \_T_1883_reg[0] ;
  wire \_T_1883_reg[1] ;
  wire _T_1927;
  wire [12:0]_T_200__0;
  wire [0:0]_T_216;
  wire _T_217;
  wire [24:0]_T_2177;
  wire _T_2222;
  wire _T_2269;
  wire _T_2305;
  wire _T_2373;
  wire _T_2377;
  wire [24:24]_T_2518;
  wire [31:1]_T_2547;
  wire \_T_2547[15]_i_3_n_0 ;
  wire \_T_2547[23]_i_3_n_0 ;
  wire \_T_2547[28]_i_3_n_0 ;
  wire \_T_2547[29]_i_3_n_0 ;
  wire \_T_2547[30]_i_3_n_0 ;
  wire \_T_2547[31]_i_4_n_0 ;
  wire \_T_2547[31]_i_5_n_0 ;
  wire \_T_2547[31]_i_6_n_0 ;
  wire \_T_2547[7]_i_3_n_0 ;
  wire [0:0]\_T_2547_reg[16]_0 ;
  wire \_T_2547_reg[16]_1 ;
  wire \_T_2547_reg[1]_0 ;
  wire [4:0]\_T_2547_reg[31]_0 ;
  wire [31:1]_T_2549;
  wire [20:1]_T_2770;
  wire [0:0]\_T_281_reg[0] ;
  wire [0:0]\_T_281_reg[3] ;
  wire \_T_294_reg[0] ;
  wire \_T_294_reg[0]_0 ;
  wire [0:0]\_T_294_reg[0]_1 ;
  wire \_T_294_reg[3] ;
  wire [0:0]_T_382;
  wire [0:0]_T_382_0;
  wire [2:0]_T_382__0;
  wire [0:0]\_T_389_reg[7] ;
  wire _T_4068_ae_ld_reg;
  wire _T_4068_pf_ld_reg;
  wire _T_4068_pf_ld_reg_0;
  wire _T_4068_pf_ld_reg_1;
  wire _T_4068_pf_ld_reg_2;
  wire _T_4068_pf_ld_reg_3;
  wire _T_4068_pf_st_reg;
  wire _T_4068_pf_st_reg_0;
  wire _T_4068_pf_st_reg_1;
  wire [0:0]_T_480;
  wire _T_481;
  wire [34:0]_T_4899;
  wire [5:0]_T_5044;
  wire _T_5074;
  wire [0:0]_T_726;
  wire [0:0]_T_877;
  wire [14:0]_T_889;
  wire [4:0]_T_909;
  wire _T_931;
  wire \_T_973_reg[1] ;
  wire [63:0]\a_data_reg[63] ;
  wire \alu/_T_198 ;
  wire \alu/_T_205 ;
  wire [7:6]\alu/_T_206 ;
  wire \alu/_T_32 ;
  wire \alu/_T_55 ;
  wire [62:0]\alu/shin ;
  wire alu_io_cmp_out;
  wire [62:0]alu_io_in1;
  wire [62:0]alu_io_in2;
  wire [32:0]alu_io_out;
  wire bad_va;
  wire [3:3]\bpu/_GEN_6 ;
  wire \buf__data_reg[12] ;
  wire \buf__data_reg[1] ;
  wire \buf__data_reg[1]_0 ;
  wire \buf__data_reg[1]_1 ;
  wire \buf__data_reg[1]_2 ;
  wire [1:0]\buf__data_reg[1]_3 ;
  wire \buf__data_reg[2] ;
  wire \buf__data_reg[3] ;
  wire \buf__data_reg[3]_0 ;
  wire [3:0]\buf__data_reg[3]_1 ;
  wire [1:0]\buf__data_reg[3]_2 ;
  wire [3:0]\buf__data_reg[3]_3 ;
  wire \buf__data_reg[4] ;
  wire \buf__data_reg[4]_0 ;
  wire buf__pc;
  wire buf__replay;
  wire buf__xcpt_ae_inst;
  wire buf__xcpt_pf_inst_reg;
  wire buf__xcpt_pf_inst_reg_0;
  wire buf__xcpt_pf_inst_reg_1;
  wire buf__xcpt_pf_inst_reg_2;
  wire \bypass_mux_1[0]_i_2_n_0 ;
  wire \bypass_mux_1[0]_i_3_n_0 ;
  wire \bypass_mux_1[0]_i_4_n_0 ;
  wire \bypass_mux_1[0]_i_5_n_0 ;
  wire \bypass_mux_1[0]_i_6_n_0 ;
  wire \bypass_mux_1[10]_i_2_n_0 ;
  wire \bypass_mux_1[10]_i_3_n_0 ;
  wire \bypass_mux_1[10]_i_4_n_0 ;
  wire \bypass_mux_1[11]_i_3_n_0 ;
  wire \bypass_mux_1[11]_i_4_n_0 ;
  wire \bypass_mux_1[11]_i_5_n_0 ;
  wire \bypass_mux_1[12]_i_2_n_0 ;
  wire \bypass_mux_1[12]_i_3_n_0 ;
  wire \bypass_mux_1[12]_i_4_n_0 ;
  wire \bypass_mux_1[13]_i_2_n_0 ;
  wire \bypass_mux_1[13]_i_3_n_0 ;
  wire \bypass_mux_1[13]_i_4_n_0 ;
  wire \bypass_mux_1[14]_i_2_n_0 ;
  wire \bypass_mux_1[14]_i_3_n_0 ;
  wire \bypass_mux_1[14]_i_4_n_0 ;
  wire \bypass_mux_1[15]_i_3_n_0 ;
  wire \bypass_mux_1[15]_i_4_n_0 ;
  wire \bypass_mux_1[15]_i_5_n_0 ;
  wire \bypass_mux_1[16]_i_2_n_0 ;
  wire \bypass_mux_1[16]_i_3_n_0 ;
  wire \bypass_mux_1[16]_i_4_n_0 ;
  wire \bypass_mux_1[17]_i_2_n_0 ;
  wire \bypass_mux_1[17]_i_3_n_0 ;
  wire \bypass_mux_1[17]_i_4_n_0 ;
  wire \bypass_mux_1[18]_i_2_n_0 ;
  wire \bypass_mux_1[18]_i_3_n_0 ;
  wire \bypass_mux_1[18]_i_4_n_0 ;
  wire \bypass_mux_1[19]_i_3_n_0 ;
  wire \bypass_mux_1[19]_i_4_n_0 ;
  wire \bypass_mux_1[19]_i_5_n_0 ;
  wire \bypass_mux_1[1]_i_2_n_0 ;
  wire \bypass_mux_1[1]_i_3_n_0 ;
  wire \bypass_mux_1[1]_i_4_n_0 ;
  wire \bypass_mux_1[1]_i_5_n_0 ;
  wire \bypass_mux_1[20]_i_2_n_0 ;
  wire \bypass_mux_1[20]_i_3_n_0 ;
  wire \bypass_mux_1[20]_i_4_n_0 ;
  wire \bypass_mux_1[21]_i_2_n_0 ;
  wire \bypass_mux_1[21]_i_3_n_0 ;
  wire \bypass_mux_1[21]_i_4_n_0 ;
  wire \bypass_mux_1[22]_i_2_n_0 ;
  wire \bypass_mux_1[22]_i_3_n_0 ;
  wire \bypass_mux_1[22]_i_4_n_0 ;
  wire \bypass_mux_1[23]_i_3_n_0 ;
  wire \bypass_mux_1[23]_i_4_n_0 ;
  wire \bypass_mux_1[23]_i_5_n_0 ;
  wire \bypass_mux_1[24]_i_2_n_0 ;
  wire \bypass_mux_1[24]_i_3_n_0 ;
  wire \bypass_mux_1[24]_i_4_n_0 ;
  wire \bypass_mux_1[25]_i_2_n_0 ;
  wire \bypass_mux_1[25]_i_3_n_0 ;
  wire \bypass_mux_1[25]_i_4_n_0 ;
  wire \bypass_mux_1[26]_i_2_n_0 ;
  wire \bypass_mux_1[26]_i_3_n_0 ;
  wire \bypass_mux_1[26]_i_4_n_0 ;
  wire \bypass_mux_1[27]_i_3_n_0 ;
  wire \bypass_mux_1[27]_i_4_n_0 ;
  wire \bypass_mux_1[27]_i_5_n_0 ;
  wire \bypass_mux_1[28]_i_2_n_0 ;
  wire \bypass_mux_1[28]_i_3_n_0 ;
  wire \bypass_mux_1[28]_i_4_n_0 ;
  wire \bypass_mux_1[29]_i_2_n_0 ;
  wire \bypass_mux_1[29]_i_3_n_0 ;
  wire \bypass_mux_1[29]_i_4_n_0 ;
  wire \bypass_mux_1[2]_i_2_n_0 ;
  wire \bypass_mux_1[2]_i_3_n_0 ;
  wire \bypass_mux_1[2]_i_4_n_0 ;
  wire \bypass_mux_1[30]_i_2_n_0 ;
  wire \bypass_mux_1[30]_i_3_n_0 ;
  wire \bypass_mux_1[30]_i_4_n_0 ;
  wire \bypass_mux_1[32]_i_2_n_0 ;
  wire \bypass_mux_1[32]_i_3_n_0 ;
  wire \bypass_mux_1[32]_i_4_n_0 ;
  wire \bypass_mux_1[3]_i_3_n_0 ;
  wire \bypass_mux_1[3]_i_4_n_0 ;
  wire \bypass_mux_1[3]_i_5_n_0 ;
  wire \bypass_mux_1[4]_i_2_n_0 ;
  wire \bypass_mux_1[4]_i_3_n_0 ;
  wire \bypass_mux_1[4]_i_4_n_0 ;
  wire \bypass_mux_1[5]_i_2_n_0 ;
  wire \bypass_mux_1[5]_i_3_n_0 ;
  wire \bypass_mux_1[5]_i_4_n_0 ;
  wire \bypass_mux_1[6]_i_2_n_0 ;
  wire \bypass_mux_1[6]_i_4_n_0 ;
  wire \bypass_mux_1[7]_i_3_n_0 ;
  wire \bypass_mux_1[7]_i_6_n_0 ;
  wire \bypass_mux_1[8]_i_2_n_0 ;
  wire \bypass_mux_1[8]_i_3_n_0 ;
  wire \bypass_mux_1[8]_i_4_n_0 ;
  wire \bypass_mux_1[9]_i_2_n_0 ;
  wire \bypass_mux_1[9]_i_3_n_0 ;
  wire \bypass_mux_1[9]_i_4_n_0 ;
  wire \bypass_mux_1_reg[0]_0 ;
  wire \bypass_mux_1_reg[17]_0 ;
  wire \bypass_mux_1_reg[18]_0 ;
  wire \bypass_mux_1_reg[19]_0 ;
  wire [3:0]\bypass_mux_1_reg[1]_0 ;
  wire \bypass_mux_1_reg[1]_1 ;
  wire \bypass_mux_1_reg[1]_2 ;
  wire \bypass_mux_1_reg[20]_0 ;
  wire \bypass_mux_1_reg[21]_0 ;
  wire \bypass_mux_1_reg[22]_0 ;
  wire \bypass_mux_1_reg[23]_0 ;
  wire \bypass_mux_1_reg[29]_0 ;
  wire \bypass_mux_1_reg[29]_1 ;
  wire \bypass_mux_1_reg[29]_2 ;
  wire \bypass_mux_1_reg[29]_3 ;
  wire \bypass_mux_1_reg[29]_4 ;
  wire \bypass_mux_1_reg[2]_0 ;
  wire \bypass_mux_1_reg[32]_0 ;
  wire \bypass_mux_1_reg[33]_0 ;
  wire \bypass_mux_1_reg[33]_1 ;
  wire \bypass_mux_1_reg[33]_2 ;
  wire \bypass_mux_1_reg[33]_3 ;
  wire \bypass_mux_1_reg[33]_4 ;
  wire \bypass_mux_1_reg[34]_0 ;
  wire \bypass_mux_1_reg[34]_1 ;
  wire \bypass_mux_1_reg[34]_2 ;
  wire \bypass_mux_1_reg[34]_3 ;
  wire \bypass_mux_1_reg[34]_4 ;
  wire \bypass_mux_1_reg[35]_0 ;
  wire \bypass_mux_1_reg[35]_1 ;
  wire \bypass_mux_1_reg[35]_2 ;
  wire \bypass_mux_1_reg[35]_3 ;
  wire \bypass_mux_1_reg[36]_0 ;
  wire \bypass_mux_1_reg[36]_1 ;
  wire [0:0]\bypass_mux_1_reg[36]_2 ;
  wire \bypass_mux_1_reg[37]_0 ;
  wire \bypass_mux_1_reg[37]_1 ;
  wire \bypass_mux_1_reg[37]_2 ;
  wire \bypass_mux_1_reg[38]_0 ;
  wire \bypass_mux_1_reg[38]_1 ;
  wire \bypass_mux_1_reg[38]_2 ;
  wire [0:0]\bypass_mux_1_reg[38]_3 ;
  wire \bypass_mux_1_reg[39]_0 ;
  wire \bypass_mux_1_reg[39]_1 ;
  wire \bypass_mux_1_reg[39]_2 ;
  wire \bypass_mux_1_reg[3]_0 ;
  wire \bypass_mux_1_reg[40]_0 ;
  wire \bypass_mux_1_reg[40]_1 ;
  wire \bypass_mux_1_reg[40]_2 ;
  wire \bypass_mux_1_reg[41]_0 ;
  wire \bypass_mux_1_reg[41]_1 ;
  wire \bypass_mux_1_reg[41]_2 ;
  wire \bypass_mux_1_reg[42]_0 ;
  wire \bypass_mux_1_reg[42]_1 ;
  wire \bypass_mux_1_reg[42]_2 ;
  wire \bypass_mux_1_reg[43]_0 ;
  wire \bypass_mux_1_reg[43]_1 ;
  wire \bypass_mux_1_reg[43]_2 ;
  wire \bypass_mux_1_reg[44]_0 ;
  wire \bypass_mux_1_reg[44]_1 ;
  wire \bypass_mux_1_reg[44]_2 ;
  wire \bypass_mux_1_reg[45]_0 ;
  wire \bypass_mux_1_reg[45]_1 ;
  wire \bypass_mux_1_reg[45]_2 ;
  wire \bypass_mux_1_reg[46]_0 ;
  wire \bypass_mux_1_reg[46]_1 ;
  wire \bypass_mux_1_reg[46]_2 ;
  wire \bypass_mux_1_reg[47]_0 ;
  wire \bypass_mux_1_reg[47]_1 ;
  wire \bypass_mux_1_reg[47]_2 ;
  wire \bypass_mux_1_reg[48]_0 ;
  wire \bypass_mux_1_reg[48]_1 ;
  wire \bypass_mux_1_reg[48]_2 ;
  wire \bypass_mux_1_reg[48]_3 ;
  wire \bypass_mux_1_reg[49]_0 ;
  wire \bypass_mux_1_reg[49]_1 ;
  wire \bypass_mux_1_reg[49]_2 ;
  wire \bypass_mux_1_reg[4]_0 ;
  wire \bypass_mux_1_reg[50]_0 ;
  wire \bypass_mux_1_reg[50]_1 ;
  wire \bypass_mux_1_reg[50]_2 ;
  wire \bypass_mux_1_reg[50]_3 ;
  wire \bypass_mux_1_reg[51]_0 ;
  wire \bypass_mux_1_reg[51]_1 ;
  wire \bypass_mux_1_reg[51]_2 ;
  wire \bypass_mux_1_reg[51]_3 ;
  wire \bypass_mux_1_reg[52]_0 ;
  wire \bypass_mux_1_reg[52]_1 ;
  wire \bypass_mux_1_reg[52]_2 ;
  wire \bypass_mux_1_reg[52]_3 ;
  wire \bypass_mux_1_reg[53]_0 ;
  wire \bypass_mux_1_reg[53]_1 ;
  wire \bypass_mux_1_reg[53]_2 ;
  wire \bypass_mux_1_reg[53]_3 ;
  wire \bypass_mux_1_reg[54]_0 ;
  wire \bypass_mux_1_reg[54]_1 ;
  wire \bypass_mux_1_reg[54]_2 ;
  wire \bypass_mux_1_reg[54]_3 ;
  wire \bypass_mux_1_reg[55]_0 ;
  wire \bypass_mux_1_reg[55]_1 ;
  wire \bypass_mux_1_reg[55]_2 ;
  wire \bypass_mux_1_reg[55]_3 ;
  wire \bypass_mux_1_reg[56]_0 ;
  wire \bypass_mux_1_reg[56]_1 ;
  wire \bypass_mux_1_reg[56]_2 ;
  wire \bypass_mux_1_reg[56]_3 ;
  wire \bypass_mux_1_reg[57]_0 ;
  wire \bypass_mux_1_reg[57]_1 ;
  wire \bypass_mux_1_reg[57]_2 ;
  wire \bypass_mux_1_reg[57]_3 ;
  wire \bypass_mux_1_reg[58]_0 ;
  wire \bypass_mux_1_reg[58]_1 ;
  wire \bypass_mux_1_reg[58]_2 ;
  wire \bypass_mux_1_reg[58]_3 ;
  wire \bypass_mux_1_reg[59]_0 ;
  wire \bypass_mux_1_reg[59]_1 ;
  wire \bypass_mux_1_reg[59]_2 ;
  wire \bypass_mux_1_reg[59]_3 ;
  wire \bypass_mux_1_reg[60]_0 ;
  wire \bypass_mux_1_reg[60]_1 ;
  wire \bypass_mux_1_reg[61]_0 ;
  wire \bypass_mux_1_reg[61]_1 ;
  wire \bypass_mux_1_reg[62]_0 ;
  wire \bypass_mux_1_reg[62]_1 ;
  wire \bypass_mux_1_reg[63]_0 ;
  wire [0:0]\bypass_mux_1_reg[63]_1 ;
  wire [0:0]\bypass_mux_1_reg[63]_2 ;
  wire \bypass_mux_1_reg[6]_0 ;
  wire [2:0]\bypass_mux_1_reg[6]_1 ;
  wire \bypass_mux_1_reg_n_0_[0] ;
  wire \bypass_mux_1_reg_n_0_[10] ;
  wire \bypass_mux_1_reg_n_0_[11] ;
  wire \bypass_mux_1_reg_n_0_[12] ;
  wire \bypass_mux_1_reg_n_0_[13] ;
  wire \bypass_mux_1_reg_n_0_[14] ;
  wire \bypass_mux_1_reg_n_0_[15] ;
  wire \bypass_mux_1_reg_n_0_[16] ;
  wire \bypass_mux_1_reg_n_0_[17] ;
  wire \bypass_mux_1_reg_n_0_[18] ;
  wire \bypass_mux_1_reg_n_0_[19] ;
  wire \bypass_mux_1_reg_n_0_[20] ;
  wire \bypass_mux_1_reg_n_0_[21] ;
  wire \bypass_mux_1_reg_n_0_[22] ;
  wire \bypass_mux_1_reg_n_0_[23] ;
  wire \bypass_mux_1_reg_n_0_[24] ;
  wire \bypass_mux_1_reg_n_0_[25] ;
  wire \bypass_mux_1_reg_n_0_[26] ;
  wire \bypass_mux_1_reg_n_0_[27] ;
  wire \bypass_mux_1_reg_n_0_[28] ;
  wire \bypass_mux_1_reg_n_0_[29] ;
  wire \bypass_mux_1_reg_n_0_[2] ;
  wire \bypass_mux_1_reg_n_0_[30] ;
  wire \bypass_mux_1_reg_n_0_[31] ;
  wire \bypass_mux_1_reg_n_0_[32] ;
  wire \bypass_mux_1_reg_n_0_[33] ;
  wire \bypass_mux_1_reg_n_0_[34] ;
  wire \bypass_mux_1_reg_n_0_[35] ;
  wire \bypass_mux_1_reg_n_0_[36] ;
  wire \bypass_mux_1_reg_n_0_[37] ;
  wire \bypass_mux_1_reg_n_0_[4] ;
  wire \bypass_mux_1_reg_n_0_[5] ;
  wire \bypass_mux_1_reg_n_0_[6] ;
  wire \bypass_mux_1_reg_n_0_[7] ;
  wire \bypass_mux_1_reg_n_0_[8] ;
  wire \bypass_mux_1_reg_n_0_[9] ;
  wire [3:0]\bypass_mux_2_reg[31]_0 ;
  wire \bypass_mux_2_reg[35]_0 ;
  wire \bypass_mux_2_reg[38]_0 ;
  wire [0:0]\bypass_mux_2_reg[63]_0 ;
  wire [0:0]\bypass_mux_2_reg[63]_1 ;
  wire [61:0]\bypass_mux_2_reg[63]_2 ;
  wire [0:0]\bypass_mux_2_reg[9]_0 ;
  wire core__115_i_2_n_0;
  wire core__116_i_10_n_0;
  wire core__116_i_11_n_0;
  wire core__130_i_5_n_0;
  wire core__131_i_3_n_0;
  wire core__131_i_4_n_0;
  wire core__131_i_5_n_0;
  wire core__132_i_3_n_0;
  wire core__132_i_4_n_0;
  wire core__132_i_5_n_0;
  wire core__133_i_4_n_0;
  wire core__133_i_5_n_0;
  wire core__133_i_6_n_0;
  wire core__134_i_10_n_0;
  wire core__134_i_11_n_0;
  wire core__134_i_3_n_0;
  wire core__134_i_4_n_0;
  wire core__134_i_5_n_0;
  wire core__134_i_6_n_0;
  wire core__134_i_7_n_0;
  wire core__134_i_8_n_0;
  wire core__134_i_9_n_0;
  wire core__135_i_10_n_0;
  wire core__135_i_11_n_0;
  wire core__135_i_3_n_0;
  wire core__135_i_4_n_0;
  wire core__135_i_5_n_0;
  wire core__135_i_6_n_0;
  wire core__135_i_7_n_0;
  wire core__135_i_8_n_0;
  wire core__135_i_9_n_0;
  wire core__136_i_10_n_0;
  wire core__136_i_11_n_0;
  wire core__136_i_3_n_0;
  wire core__136_i_4_n_0;
  wire core__136_i_5_n_0;
  wire core__136_i_6_n_0;
  wire core__136_i_7_n_0;
  wire core__136_i_8_n_0;
  wire core__136_i_9_n_0;
  wire core__137_i_10_n_0;
  wire core__137_i_11_n_0;
  wire core__137_i_4_n_0;
  wire core__137_i_5_n_0;
  wire core__137_i_6_n_0;
  wire core__137_i_7_n_0;
  wire core__137_i_8_n_0;
  wire core__137_i_9_n_0;
  wire core__138_i_3_n_0;
  wire core__138_i_4_n_0;
  wire core__138_i_5_n_0;
  wire core__138_i_6_n_0;
  wire core__138_i_7_n_0;
  wire core__138_i_8_n_0;
  wire core__139_i_3_n_0;
  wire core__139_i_4_n_0;
  wire core__139_i_5_n_0;
  wire core__139_i_6_n_0;
  wire core__139_i_7_n_0;
  wire core__139_i_8_n_0;
  wire core__140_i_10_n_0;
  wire core__140_i_3_n_0;
  wire core__140_i_4_n_0;
  wire core__140_i_5_n_0;
  wire core__140_i_6_n_0;
  wire core__140_i_7_n_0;
  wire core__140_i_8_n_0;
  wire core__140_i_9_n_0;
  wire core__141_i_10_n_0;
  wire core__141_i_4_n_0;
  wire core__141_i_5_n_0;
  wire core__141_i_6_n_0;
  wire core__141_i_7_n_0;
  wire core__141_i_8_n_0;
  wire core__141_i_9_n_0;
  wire core__142_i_3_n_0;
  wire core__142_i_4_n_0;
  wire core__142_i_5_n_0;
  wire core__142_i_6_n_0;
  wire core__142_i_7_n_0;
  wire core__142_i_8_n_0;
  wire core__142_i_9_n_0;
  wire core__143_i_3_n_0;
  wire core__143_i_4_n_0;
  wire core__143_i_5_n_0;
  wire core__143_i_6_n_0;
  wire core__143_i_7_n_0;
  wire core__144_i_3_n_0;
  wire core__144_i_4_n_0;
  wire core__144_i_5_n_0;
  wire core__144_i_6_n_0;
  wire core__144_i_7_n_0;
  wire core__144_i_8_n_0;
  wire core__145_i_5_n_0;
  wire core__145_i_7_n_0;
  wire core__146_i_4_n_0;
  wire core__146_i_5_n_0;
  wire core__146_i_6_n_0;
  wire core__147_i_4_n_0;
  wire core__147_i_5_n_0;
  wire core__147_i_6_n_0;
  wire core__148_i_4_n_0;
  wire core__148_i_5_n_0;
  wire core__148_i_6_n_0;
  wire core__149_i_5_n_0;
  wire core__149_i_6_n_0;
  wire core__149_i_7_n_0;
  wire core__150_i_4_n_0;
  wire core__150_i_5_n_0;
  wire core__150_i_6_n_0;
  wire core__151_i_4_n_0;
  wire core__151_i_5_n_0;
  wire core__151_i_6_n_0;
  wire core__152_i_4_n_0;
  wire core__152_i_5_n_0;
  wire core__152_i_6_n_0;
  wire core__153_i_5_n_0;
  wire core__153_i_6_n_0;
  wire core__153_i_7_n_0;
  wire core__154_i_10_n_0;
  wire core__154_i_11_n_0;
  wire core__154_i_12_n_0;
  wire core__154_i_4_n_0;
  wire core__154_i_5_n_0;
  wire core__154_i_6_n_0;
  wire core__154_i_7_n_0;
  wire core__154_i_8_n_0;
  wire core__154_i_9_n_0;
  wire core__155_i_4_n_0;
  wire core__155_i_5_n_0;
  wire core__155_i_6_n_0;
  wire core__156_i_4_n_0;
  wire core__156_i_5_n_0;
  wire core__156_i_6_n_0;
  wire core__157_i_4_n_0;
  wire core__157_i_5_n_0;
  wire core__157_i_6_n_0;
  wire core__157_i_7_n_0;
  wire core__158_i_3_n_0;
  wire core__158_i_4_n_0;
  wire core__158_i_5_n_0;
  wire core__158_i_6_n_0;
  wire core__158_i_7_n_0;
  wire core__159_i_10_n_0;
  wire core__159_i_11_n_0;
  wire core__159_i_12_n_0;
  wire core__159_i_13_n_0;
  wire core__159_i_14_n_0;
  wire core__159_i_15_n_0;
  wire core__159_i_3_n_0;
  wire core__159_i_4_n_0;
  wire core__159_i_5_n_0;
  wire core__159_i_6_n_0;
  wire core__159_i_7_n_0;
  wire core__159_i_8_n_0;
  wire core__159_i_9_n_0;
  wire core__160_i_2_n_0;
  wire core__160_i_3_n_0;
  wire core__160_i_4_n_0;
  wire core__160_i_5_n_0;
  wire core__160_i_6_n_0;
  wire core__160_i_7_n_0;
  wire core__160_i_8_n_0;
  wire core__161_i_3_n_0;
  wire core__161_i_4_n_0;
  wire core__161_i_5_n_0;
  wire core__161_i_6_n_0;
  wire core__162_i_5_n_0;
  wire core__162_i_6_n_0;
  wire core__163_i_5_n_0;
  wire core__163_i_6_n_0;
  wire core__163_i_7_n_0;
  wire core__163_i_8_n_0;
  wire core__166_i_5_n_0;
  wire core__166_i_6_n_0;
  wire core__168_i_5_n_0;
  wire core__436_i_3_n_0;
  wire core__441_i_3_n_0;
  wire core__506_i_2_n_0;
  wire core__638_i_4_n_0;
  wire core__639_i_10_n_0;
  wire core__639_i_11_n_0;
  wire core__641_i_12_n_0;
  wire core__641_i_13_n_0;
  wire core__643_i_12_n_0;
  wire core__643_i_13_n_0;
  wire core__644_i_12_n_0;
  wire core__644_i_13_n_0;
  wire core__649_i_10_n_0;
  wire core__649_i_11_n_0;
  wire core__649_i_12_n_0;
  wire core__649_i_5_n_0;
  wire core__649_i_6_n_0;
  wire core__649_i_7_n_0;
  wire core__649_i_8_n_0;
  wire core__649_i_9_n_0;
  wire core__650_i_2_n_0;
  wire core__651_i_2_n_0;
  wire core__652_i_2_n_0;
  wire core__653_i_2_n_0;
  wire core__654_i_2_n_0;
  wire core__655_i_2_n_0;
  wire core__656_i_2_n_0;
  wire core__657_i_2_n_0;
  wire core__658_i_2_n_0;
  wire core__707_i_3_n_0;
  wire core__707_i_4_n_0;
  wire \count_reg[0] ;
  wire \count_reg[1] ;
  wire \count_reg[1]_0 ;
  wire \count_reg[1]_1 ;
  wire \count_reg[1]_2 ;
  wire [37:4]csr_io_bp_0_address;
  wire csr_io_bp_0_control_action;
  wire csr_io_bp_0_control_m;
  wire csr_io_bp_0_control_s;
  wire csr_io_bp_0_control_u;
  wire csr_io_interrupt;
  wire [8:3]csr_io_rw_addr;
  wire csr_io_status_debug;
  wire [0:0]csr_io_tval;
  wire csr_n_636;
  wire csr_n_637;
  wire csr_n_638;
  wire csr_n_639;
  wire csr_n_641;
  wire csr_n_642;
  wire csr_n_643;
  wire csr_n_644;
  wire csr_n_664;
  wire csr_n_665;
  wire csr_n_666;
  wire csr_n_667;
  wire csr_n_668;
  wire csr_n_669;
  wire csr_n_670;
  wire csr_n_671;
  wire csr_n_672;
  wire csr_n_673;
  wire csr_n_674;
  wire csr_n_675;
  wire csr_n_676;
  wire csr_n_677;
  wire csr_n_678;
  wire csr_n_679;
  wire csr_n_680;
  wire csr_n_681;
  wire csr_n_682;
  wire csr_n_683;
  wire csr_n_684;
  wire csr_n_685;
  wire csr_n_686;
  wire csr_n_687;
  wire csr_n_688;
  wire csr_n_689;
  wire csr_n_690;
  wire csr_n_691;
  wire csr_n_692;
  wire csr_n_693;
  wire csr_n_694;
  wire csr_n_695;
  wire csr_n_696;
  wire csr_n_697;
  wire csr_n_698;
  wire csr_n_699;
  wire csr_n_700;
  wire csr_n_701;
  wire csr_n_702;
  wire csr_n_703;
  wire csr_n_747;
  wire csr_n_748;
  wire data_arrays_0_0_reg_i_53_n_0;
  wire dcacheArb_io_requestor_1_ordered;
  wire dcacheArb_io_requestor_1_replay_next;
  wire [32:0]dcacheArb_io_requestor_1_req_bits_addr;
  wire [2:0]dcacheArb_io_requestor_1_req_bits_typ;
  wire dcacheArb_io_requestor_1_req_ready;
  wire dcacheArb_io_requestor_1_req_valid;
  wire [43:0]dcacheArb_io_requestor_1_resp_bits_data;
  wire [63:0]dcacheArb_io_requestor_1_resp_bits_data_word_bypass;
  wire dcacheArb_io_requestor_1_resp_bits_replay;
  wire dcacheArb_io_requestor_1_resp_valid;
  wire dcacheArb_io_requestor_1_s1_kill;
  wire dcacheArb_io_requestor_1_s2_nack;
  wire dcacheArb_io_requestor_1_s2_xcpt_ma_ld;
  wire dcacheArb_io_requestor_1_s2_xcpt_ma_st;
  wire dcacheArb_io_requestor_1_s2_xcpt_pf_ld;
  wire dcacheArb_io_requestor_1_s2_xcpt_pf_st;
  wire dcache_blocked;
  wire dcache_blocked0;
  wire dcache_io_cpu_invalidate_lr;
  wire dcache_io_ptw_resp_bits_ae;
  wire dcache_io_ptw_resp_bits_homogeneous;
  wire [1:0]dcache_io_ptw_resp_bits_level;
  wire dcache_io_ptw_resp_valid;
  wire dcache_io_ptw_status_mxr;
  wire dcache_io_ptw_status_sum;
  wire div_n_138;
  wire div_n_139;
  wire div_n_140;
  wire div_n_141;
  wire div_n_142;
  wire div_n_143;
  wire div_n_144;
  wire div_n_145;
  wire div_n_146;
  wire div_n_147;
  wire div_n_148;
  wire div_n_149;
  wire div_n_150;
  wire div_n_151;
  wire div_n_152;
  wire div_n_153;
  wire div_n_154;
  wire div_n_155;
  wire div_n_156;
  wire div_n_157;
  wire div_n_158;
  wire div_n_159;
  wire div_n_160;
  wire div_n_161;
  wire div_n_162;
  wire div_n_163;
  wire div_n_164;
  wire div_n_165;
  wire div_n_166;
  wire div_n_167;
  wire div_n_170;
  wire div_n_218;
  wire div_n_219;
  wire div_n_220;
  wire div_n_221;
  wire div_n_222;
  wire div_n_223;
  wire div_n_224;
  wire div_n_225;
  wire div_n_226;
  wire div_n_227;
  wire div_n_228;
  wire div_n_229;
  wire div_n_230;
  wire div_n_234;
  wire div_n_235;
  wire div_n_236;
  wire div_n_237;
  wire div_n_238;
  wire div_n_239;
  wire div_n_240;
  wire div_n_368;
  wire div_n_526;
  wire [2:0]\divisor_reg[15] ;
  wire [3:0]\divisor_reg[15]_0 ;
  wire [3:0]\divisor_reg[15]_1 ;
  wire [3:0]\divisor_reg[15]_2 ;
  wire [3:0]\divisor_reg[15]_3 ;
  wire [3:0]\divisor_reg[15]_4 ;
  wire [3:0]\divisor_reg[15]_5 ;
  wire [3:0]\divisor_reg[15]_6 ;
  wire [3:0]\divisor_reg[15]_7 ;
  wire [1:0]\divisor_reg[15]_8 ;
  wire [0:0]\divisor_reg[18] ;
  wire [0:0]\divisor_reg[1] ;
  wire [2:0]\divisor_reg[32] ;
  wire [3:0]\divisor_reg[32]_0 ;
  wire [3:0]\divisor_reg[32]_1 ;
  wire [0:0]\divisor_reg[35] ;
  wire [3:0]\divisor_reg[51] ;
  wire [0:0]\divisor_reg[52] ;
  wire [5:0]\divisor_reg[57] ;
  wire doUncachedResp_reg;
  wire [15:0]\elts_0_data_reg[15] ;
  wire [0:0]\elts_0_pc_reg[38] ;
  wire [18:0]\elts_0_pc_reg[39] ;
  wire elts_0_xcpt_ae_inst_reg;
  wire [63:0]ex_cause;
  wire [0:0]\ex_cause_reg[1]_0 ;
  wire [0:0]\ex_cause_reg[1]_1 ;
  wire [3:0]\ex_cause_reg[1]_10 ;
  wire [3:0]\ex_cause_reg[1]_11 ;
  wire [3:0]\ex_cause_reg[1]_12 ;
  wire [2:0]\ex_cause_reg[1]_13 ;
  wire [2:0]\ex_cause_reg[1]_14 ;
  wire [2:0]\ex_cause_reg[1]_2 ;
  wire [2:0]\ex_cause_reg[1]_3 ;
  wire [3:0]\ex_cause_reg[1]_4 ;
  wire [3:0]\ex_cause_reg[1]_5 ;
  wire [3:0]\ex_cause_reg[1]_6 ;
  wire [3:0]\ex_cause_reg[1]_7 ;
  wire [3:0]\ex_cause_reg[1]_8 ;
  wire [3:0]\ex_cause_reg[1]_9 ;
  wire ex_ctrl_alu_dw_reg_0;
  wire ex_ctrl_alu_dw_reg_1;
  wire ex_ctrl_alu_dw_reg_10;
  wire ex_ctrl_alu_dw_reg_11;
  wire ex_ctrl_alu_dw_reg_12;
  wire ex_ctrl_alu_dw_reg_13;
  wire ex_ctrl_alu_dw_reg_14;
  wire ex_ctrl_alu_dw_reg_15;
  wire ex_ctrl_alu_dw_reg_16;
  wire ex_ctrl_alu_dw_reg_17;
  wire ex_ctrl_alu_dw_reg_18;
  wire ex_ctrl_alu_dw_reg_19;
  wire ex_ctrl_alu_dw_reg_2;
  wire ex_ctrl_alu_dw_reg_20;
  wire ex_ctrl_alu_dw_reg_21;
  wire ex_ctrl_alu_dw_reg_22;
  wire ex_ctrl_alu_dw_reg_23;
  wire ex_ctrl_alu_dw_reg_24;
  wire ex_ctrl_alu_dw_reg_25;
  wire ex_ctrl_alu_dw_reg_26;
  wire ex_ctrl_alu_dw_reg_27;
  wire ex_ctrl_alu_dw_reg_28;
  wire ex_ctrl_alu_dw_reg_29;
  wire ex_ctrl_alu_dw_reg_3;
  wire ex_ctrl_alu_dw_reg_30;
  wire ex_ctrl_alu_dw_reg_31;
  wire ex_ctrl_alu_dw_reg_32;
  wire ex_ctrl_alu_dw_reg_33;
  wire ex_ctrl_alu_dw_reg_4;
  wire ex_ctrl_alu_dw_reg_5;
  wire ex_ctrl_alu_dw_reg_6;
  wire ex_ctrl_alu_dw_reg_7;
  wire ex_ctrl_alu_dw_reg_8;
  wire ex_ctrl_alu_dw_reg_9;
  wire [2:0]ex_ctrl_alu_fn;
  wire \ex_ctrl_alu_fn_reg[3]_0 ;
  wire \ex_ctrl_alu_fn_reg[3]_1 ;
  wire \ex_ctrl_alu_fn_reg[3]_2 ;
  wire \ex_ctrl_alu_fn_reg[3]_3 ;
  wire \ex_ctrl_alu_fn_reg[3]_4 ;
  wire \ex_ctrl_alu_fn_reg[3]_5 ;
  wire \ex_ctrl_alu_fn_reg[3]_6 ;
  wire \ex_ctrl_alu_fn_reg[3]_7 ;
  wire \ex_ctrl_alu_fn_reg[3]_8 ;
  wire [0:0]\ex_ctrl_alu_fn_reg[3]_9 ;
  wire ex_ctrl_branch;
  wire \ex_ctrl_csr_reg[0]_0 ;
  wire \ex_ctrl_csr_reg[1]_0 ;
  wire \ex_ctrl_csr_reg[2]_0 ;
  wire ex_ctrl_div;
  wire ex_ctrl_div_reg_0;
  wire ex_ctrl_fence_i;
  wire ex_ctrl_jal;
  wire ex_ctrl_jalr;
  wire ex_ctrl_mem;
  wire ex_ctrl_mem_reg_0;
  wire ex_ctrl_mem_reg_1;
  wire ex_ctrl_mem_reg_10;
  wire ex_ctrl_mem_reg_11;
  wire ex_ctrl_mem_reg_2;
  wire ex_ctrl_mem_reg_3;
  wire ex_ctrl_mem_reg_4;
  wire ex_ctrl_mem_reg_5;
  wire ex_ctrl_mem_reg_6;
  wire ex_ctrl_mem_reg_7;
  wire ex_ctrl_mem_reg_8;
  wire ex_ctrl_mem_reg_9;
  wire [1:0]\ex_ctrl_mem_type_reg[0]_0 ;
  wire ex_ctrl_rxs2;
  wire \ex_ctrl_sel_alu1_reg[0]_0 ;
  wire \ex_ctrl_sel_alu1_reg[1]_0 ;
  wire [1:0]ex_ctrl_sel_alu2;
  wire \ex_ctrl_sel_alu2_reg[1]_0 ;
  wire \ex_ctrl_sel_alu2_reg[1]_1 ;
  wire \ex_ctrl_sel_alu2_reg[1]_2 ;
  wire \ex_ctrl_sel_alu2_reg[1]_3 ;
  wire \ex_ctrl_sel_alu2_reg[1]_4 ;
  wire \ex_ctrl_sel_alu2_reg[1]_5 ;
  wire \ex_ctrl_sel_imm_reg[1]_0 ;
  wire \ex_ctrl_sel_imm_reg[1]_1 ;
  wire ex_ctrl_wxd;
  wire ex_ctrl_wxd_reg_0;
  wire [1:0]ex_ctrl_wxd_reg_1;
  wire ex_reg_flush_pipe;
  wire \ex_reg_inst_reg[10]_0 ;
  wire \ex_reg_inst_reg[10]_1 ;
  wire \ex_reg_inst_reg[10]_2 ;
  wire \ex_reg_inst_reg[10]_3 ;
  wire \ex_reg_inst_reg[10]_4 ;
  wire \ex_reg_inst_reg[10]_5 ;
  wire \ex_reg_inst_reg[10]_6 ;
  wire \ex_reg_inst_reg[10]_7 ;
  wire [15:0]\ex_reg_inst_reg[11]_0 ;
  wire \ex_reg_inst_reg[26]_0 ;
  wire \ex_reg_inst_reg_n_0_[12] ;
  wire \ex_reg_inst_reg_n_0_[13] ;
  wire \ex_reg_inst_reg_n_0_[14] ;
  wire \ex_reg_inst_reg_n_0_[15] ;
  wire \ex_reg_inst_reg_n_0_[16] ;
  wire \ex_reg_inst_reg_n_0_[17] ;
  wire \ex_reg_inst_reg_n_0_[18] ;
  wire \ex_reg_inst_reg_n_0_[19] ;
  wire \ex_reg_inst_reg_n_0_[21] ;
  wire \ex_reg_inst_reg_n_0_[22] ;
  wire \ex_reg_inst_reg_n_0_[23] ;
  wire \ex_reg_inst_reg_n_0_[24] ;
  wire \ex_reg_inst_reg_n_0_[25] ;
  wire \ex_reg_inst_reg_n_0_[28] ;
  wire \ex_reg_inst_reg_n_0_[29] ;
  wire \ex_reg_inst_reg_n_0_[30] ;
  wire ex_reg_load_use;
  wire [39:1]ex_reg_pc;
  wire [19:0]\ex_reg_pc_reg[39]_0 ;
  wire [0:0]\ex_reg_pc_reg[39]_1 ;
  wire ex_reg_replay;
  wire ex_reg_replay0;
  wire ex_reg_rs_bypass_0;
  wire ex_reg_rs_bypass_0_reg_0;
  wire ex_reg_rs_bypass_0_reg_1;
  wire ex_reg_rs_bypass_1;
  wire ex_reg_rs_bypass_1_reg_0;
  wire [1:0]ex_reg_rs_lsb_0;
  wire \ex_reg_rs_lsb_0_reg[0]_0 ;
  wire \ex_reg_rs_lsb_0_reg[0]_1 ;
  wire \ex_reg_rs_lsb_0_reg[1]_0 ;
  wire \ex_reg_rs_lsb_1_reg_n_0_[0] ;
  wire \ex_reg_rs_lsb_1_reg_n_0_[1] ;
  wire \ex_reg_rs_msb_0_reg[10]_0 ;
  wire \ex_reg_rs_msb_0_reg[11]_0 ;
  wire \ex_reg_rs_msb_0_reg[12]_0 ;
  wire \ex_reg_rs_msb_0_reg[13]_0 ;
  wire \ex_reg_rs_msb_0_reg[14]_0 ;
  wire \ex_reg_rs_msb_0_reg[15]_0 ;
  wire \ex_reg_rs_msb_0_reg[16]_0 ;
  wire \ex_reg_rs_msb_0_reg[17]_0 ;
  wire \ex_reg_rs_msb_0_reg[18]_0 ;
  wire \ex_reg_rs_msb_0_reg[19]_0 ;
  wire \ex_reg_rs_msb_0_reg[20]_0 ;
  wire \ex_reg_rs_msb_0_reg[21]_0 ;
  wire \ex_reg_rs_msb_0_reg[22]_0 ;
  wire \ex_reg_rs_msb_0_reg[23]_0 ;
  wire \ex_reg_rs_msb_0_reg[24]_0 ;
  wire \ex_reg_rs_msb_0_reg[25]_0 ;
  wire \ex_reg_rs_msb_0_reg[26]_0 ;
  wire [19:0]\ex_reg_rs_msb_0_reg[27]_0 ;
  wire \ex_reg_rs_msb_0_reg[27]_1 ;
  wire \ex_reg_rs_msb_0_reg[8]_0 ;
  wire \ex_reg_rs_msb_0_reg[9]_0 ;
  wire \ex_reg_rs_msb_0_reg_n_0_[0] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[10] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[11] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[12] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[13] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[14] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[15] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[16] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[17] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[18] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[19] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[1] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[20] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[21] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[22] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[23] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[24] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[25] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[26] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[27] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[28] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[29] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[2] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[30] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[31] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[32] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[33] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[34] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[35] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[36] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[37] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[38] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[39] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[3] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[40] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[41] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[42] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[43] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[44] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[45] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[46] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[47] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[48] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[49] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[4] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[50] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[51] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[52] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[53] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[54] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[55] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[56] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[57] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[58] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[59] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[5] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[60] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[61] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[6] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[7] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[8] ;
  wire \ex_reg_rs_msb_0_reg_n_0_[9] ;
  wire [66:0]\ex_reg_rs_msb_1_reg[29]_0 ;
  wire \ex_reg_rs_msb_1_reg[61]_0 ;
  wire [2:0]\ex_reg_rs_msb_1_reg[61]_1 ;
  wire \ex_reg_rs_msb_1_reg[61]_2 ;
  wire \ex_reg_rs_msb_1_reg_n_0_[0] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[10] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[11] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[12] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[13] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[14] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[15] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[16] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[17] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[18] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[19] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[1] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[20] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[21] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[22] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[23] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[24] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[25] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[26] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[27] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[28] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[29] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[2] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[30] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[31] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[32] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[33] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[34] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[35] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[36] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[37] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[38] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[39] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[3] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[40] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[41] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[42] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[43] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[44] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[45] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[46] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[47] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[48] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[49] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[4] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[50] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[51] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[52] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[53] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[54] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[55] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[56] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[57] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[58] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[59] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[5] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[60] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[61] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[6] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[7] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[8] ;
  wire \ex_reg_rs_msb_1_reg_n_0_[9] ;
  wire ex_reg_rvc_reg_0;
  wire ex_reg_rvc_reg_1;
  wire ex_reg_rvc_reg_10;
  wire ex_reg_rvc_reg_11;
  wire ex_reg_rvc_reg_12;
  wire ex_reg_rvc_reg_13;
  wire ex_reg_rvc_reg_14;
  wire ex_reg_rvc_reg_15;
  wire ex_reg_rvc_reg_16;
  wire ex_reg_rvc_reg_2;
  wire ex_reg_rvc_reg_3;
  wire ex_reg_rvc_reg_4;
  wire ex_reg_rvc_reg_5;
  wire ex_reg_rvc_reg_6;
  wire ex_reg_rvc_reg_7;
  wire ex_reg_rvc_reg_8;
  wire ex_reg_rvc_reg_9;
  wire ex_reg_valid;
  wire ex_reg_xcpt;
  wire ex_reg_xcpt_interrupt;
  wire ex_reg_xcpt_interrupt0;
  wire ex_sfence;
  wire frontend_io_cpu_req_bits_speculative;
  wire [1:0]frontend_io_cpu_resp_bits_data;
  wire [38:0]frontend_io_cpu_resp_bits_pc;
  wire frontend_io_cpu_resp_bits_replay;
  wire frontend_io_cpu_resp_bits_xcpt_ae_inst;
  wire frontend_io_cpu_resp_bits_xcpt_pf_inst;
  wire frontend_io_cpu_resp_valid;
  wire frontend_io_cpu_sfence_bits_rs2;
  wire frontend_io_cpu_sfence_valid;
  wire [1:0]frontend_io_ptw_pmp_1_cfg_a;
  wire frontend_io_ptw_pmp_1_cfg_w;
  wire [1:0]frontend_io_ptw_pmp_2_cfg_a;
  wire [1:0]frontend_io_ptw_pmp_6_cfg_a;
  wire [1:0]frontend_io_ptw_pmp_7_cfg_a;
  wire [0:0]frontend_io_ptw_ptbr_mode;
  wire [1:0]frontend_io_ptw_status_prv;
  wire hitsVec_4;
  wire host_clk;
  wire [4:0]ibuf_io_inst_0_bits_inst_rd;
  wire [4:0]ibuf_io_inst_0_bits_inst_rs1;
  wire [4:0]ibuf_io_inst_0_bits_inst_rs2;
  wire [0:0]ibuf_io_inst_0_bits_raw;
  wire ibuf_io_inst_0_bits_xcpt0_ae_inst;
  wire [36:1]ibuf_io_pc;
  wire ibuf_n_47;
  wire ibuf_n_50;
  wire ibuf_n_52;
  wire ibuf_n_56;
  wire ibuf_n_64;
  wire ibuf_n_65;
  wire ibuf_n_68;
  wire ibuf_n_70;
  wire ibuf_n_71;
  wire ibuf_n_72;
  wire ibuf_n_73;
  wire ibuf_n_74;
  wire id_ctrl_fence_i;
  wire id_ctrl_jal;
  wire id_ctrl_mem;
  wire id_ctrl_rxs2;
  wire [1:0]id_ctrl_sel_alu1;
  wire id_ctrl_wxd;
  wire id_load_use;
  wire id_reg_fence_reg_0;
  wire invalidated;
  wire invalidated_reg;
  wire [0:0]io_mask;
  wire \lrscCount_reg[0] ;
  wire \lrscCount_reg[0]_0 ;
  wire mem_br_taken_;
  wire [0:0]mem_br_taken__reg_0;
  wire mem_ctrl_branch;
  wire mem_ctrl_branch_reg_0;
  wire [2:0]mem_ctrl_csr;
  wire mem_ctrl_div;
  wire mem_ctrl_fence_i_reg_0;
  wire mem_ctrl_fp;
  wire mem_ctrl_jal;
  wire mem_ctrl_jalr;
  wire mem_ctrl_mem;
  wire \mem_ctrl_mem_type_reg_n_0_[0] ;
  wire \mem_ctrl_mem_type_reg_n_0_[1] ;
  wire mem_ctrl_wxd;
  wire [63:0]mem_int_wdata;
  wire mem_pc_valid;
  wire [63:0]mem_reg_cause;
  wire mem_reg_flush_pipe;
  wire mem_reg_flush_pipe_reg_0;
  wire \mem_reg_inst_reg[11]_0 ;
  wire [7:0]\mem_reg_inst_reg[31]_0 ;
  wire [0:0]\mem_reg_inst_reg[9]_0 ;
  wire [0:0]\mem_reg_inst_reg[9]_1 ;
  wire mem_reg_load;
  wire [0:0]\mem_reg_pc_reg[31]_0 ;
  wire mem_reg_replay;
  wire mem_reg_replay0;
  wire mem_reg_replay_reg_0;
  wire [63:0]mem_reg_rs2;
  wire [63:8]mem_reg_rs20_in;
  wire \mem_reg_rs2[63]_i_1_n_0 ;
  wire \mem_reg_rs2_reg[0]_0 ;
  wire \mem_reg_rs2_reg[1]_0 ;
  wire \mem_reg_rs2_reg[25]_0 ;
  wire \mem_reg_rs2_reg[2]_0 ;
  wire \mem_reg_rs2_reg[3]_0 ;
  wire [1:0]\mem_reg_rs2_reg[3]_1 ;
  wire \mem_reg_rs2_reg[4]_0 ;
  wire \mem_reg_rs2_reg[5]_0 ;
  wire \mem_reg_rs2_reg[6]_0 ;
  wire \mem_reg_rs2_reg[7]_0 ;
  wire mem_reg_rvc;
  wire mem_reg_rvc_reg_0;
  wire mem_reg_sfence;
  wire mem_reg_sfence_reg_0;
  wire mem_reg_sfence_reg_1;
  wire mem_reg_sfence_reg_2;
  wire mem_reg_slow_bypass;
  wire mem_reg_slow_bypass_reg_0;
  wire mem_reg_slow_bypass_reg_1;
  wire mem_reg_store;
  wire mem_reg_valid;
  wire mem_reg_valid_reg_0;
  wire mem_reg_xcpt;
  wire mem_reg_xcpt0;
  wire mem_reg_xcpt_interrupt;
  wire mem_reg_xcpt_interrupt0;
  wire [1:0]mem_reg_xcpt_interrupt_reg_0;
  wire nBufValid_reg;
  wire nBufValid_reg_0;
  wire nBufValid_reg_1;
  wire nBufValid_reg_2;
  wire nBufValid_reg_3;
  wire nBufValid_reg_4;
  wire nBufValid_reg_5;
  wire [4:0]nBufValid_reg_6;
  wire nBufValid_reg_7;
  wire [2:0]nBufValid_reg_8;
  wire [0:0]nBufValid_reg_9;
  wire neg_out_reg;
  wire [63:0]out;
  wire [39:0]p_0_in;
  wire [4:0]p_0_in__0;
  wire p_13_in;
  wire p_2_in;
  wire p_31_in;
  wire [0:0]q_reg;
  wire \r_pte_ppn_reg[0] ;
  wire \r_pte_ppn_reg[10] ;
  wire \r_pte_ppn_reg[11] ;
  wire \r_pte_ppn_reg[12] ;
  wire \r_pte_ppn_reg[13] ;
  wire \r_pte_ppn_reg[14] ;
  wire \r_pte_ppn_reg[15] ;
  wire \r_pte_ppn_reg[16] ;
  wire \r_pte_ppn_reg[16]_0 ;
  wire \r_pte_ppn_reg[16]_1 ;
  wire \r_pte_ppn_reg[16]_2 ;
  wire \r_pte_ppn_reg[16]_3 ;
  wire \r_pte_ppn_reg[16]_4 ;
  wire \r_pte_ppn_reg[16]_5 ;
  wire \r_pte_ppn_reg[16]_6 ;
  wire \r_pte_ppn_reg[16]_7 ;
  wire \r_pte_ppn_reg[17] ;
  wire \r_pte_ppn_reg[18] ;
  wire [19:0]\r_pte_ppn_reg[19] ;
  wire [19:0]\r_pte_ppn_reg[19]_0 ;
  wire \r_pte_ppn_reg[1] ;
  wire \r_pte_ppn_reg[2] ;
  wire \r_pte_ppn_reg[3] ;
  wire \r_pte_ppn_reg[3]_0 ;
  wire \r_pte_ppn_reg[3]_1 ;
  wire \r_pte_ppn_reg[3]_2 ;
  wire \r_pte_ppn_reg[3]_3 ;
  wire \r_pte_ppn_reg[3]_4 ;
  wire \r_pte_ppn_reg[3]_5 ;
  wire \r_pte_ppn_reg[3]_6 ;
  wire \r_pte_ppn_reg[3]_7 ;
  wire \r_pte_ppn_reg[4] ;
  wire \r_pte_ppn_reg[5] ;
  wire \r_pte_ppn_reg[5]_0 ;
  wire \r_pte_ppn_reg[5]_1 ;
  wire \r_pte_ppn_reg[5]_2 ;
  wire \r_pte_ppn_reg[5]_3 ;
  wire \r_pte_ppn_reg[5]_4 ;
  wire \r_pte_ppn_reg[5]_5 ;
  wire \r_pte_ppn_reg[5]_6 ;
  wire \r_pte_ppn_reg[5]_7 ;
  wire \r_pte_ppn_reg[6] ;
  wire \r_pte_ppn_reg[7] ;
  wire \r_pte_ppn_reg[7]_0 ;
  wire \r_pte_ppn_reg[7]_1 ;
  wire \r_pte_ppn_reg[7]_2 ;
  wire \r_pte_ppn_reg[7]_3 ;
  wire \r_pte_ppn_reg[7]_4 ;
  wire \r_pte_ppn_reg[7]_5 ;
  wire \r_pte_ppn_reg[7]_6 ;
  wire \r_pte_ppn_reg[7]_7 ;
  wire \r_pte_ppn_reg[8] ;
  wire \r_pte_ppn_reg[9] ;
  wire \r_refill_waddr_reg[0] ;
  wire [1:0]\r_refill_waddr_reg[1] ;
  wire refill_valid;
  wire [0:0]\reg_bp_0_address_reg[36] ;
  wire \reg_bp_0_address_reg[3] ;
  wire reg_bp_0_control_action_reg;
  wire [13:0]\reg_bp_0_control_tmatch_reg[1] ;
  wire \reg_bp_0_control_tmatch_reg[1]_0 ;
  wire \reg_dcsr_cause_reg[0] ;
  wire \reg_dcsr_cause_reg[1] ;
  wire reg_dcsr_prv;
  wire reg_dcsr_step;
  wire reg_debug_reg;
  wire reg_debug_reg_0;
  wire reg_debug_reg_1;
  wire reg_debug_reg_2;
  wire \reg_dpc_reg[12] ;
  wire [38:0]\reg_dpc_reg[39] ;
  wire \reg_dscratch_reg[0] ;
  wire \reg_entries_0_reg[0] ;
  wire [0:0]\reg_entries_0_reg[0]_0 ;
  wire [0:0]\reg_entries_0_reg[0]_1 ;
  wire [0:0]\reg_entries_0_reg[0]_2 ;
  wire [0:0]\reg_entries_0_reg[0]_3 ;
  wire [0:0]\reg_entries_0_reg[0]_4 ;
  wire [0:0]\reg_entries_0_reg[0]_5 ;
  wire [0:0]\reg_entries_0_reg[0]_6 ;
  wire [0:0]\reg_entries_0_reg[0]_7 ;
  wire [0:0]\reg_entries_0_reg[10] ;
  wire \reg_entries_0_reg[4] ;
  wire \reg_entries_0_reg[4]_0 ;
  wire [2:0]\reg_entries_0_reg[4]_1 ;
  wire [3:0]\reg_entries_0_reg[4]_10 ;
  wire [3:0]\reg_entries_0_reg[4]_11 ;
  wire [3:0]\reg_entries_0_reg[4]_12 ;
  wire [2:0]\reg_entries_0_reg[4]_13 ;
  wire \reg_entries_0_reg[4]_14 ;
  wire \reg_entries_0_reg[4]_15 ;
  wire \reg_entries_0_reg[4]_16 ;
  wire \reg_entries_0_reg[4]_17 ;
  wire \reg_entries_0_reg[4]_18 ;
  wire \reg_entries_0_reg[4]_19 ;
  wire [2:0]\reg_entries_0_reg[4]_2 ;
  wire [3:0]\reg_entries_0_reg[4]_20 ;
  wire [3:0]\reg_entries_0_reg[4]_21 ;
  wire \reg_entries_0_reg[4]_22 ;
  wire [3:0]\reg_entries_0_reg[4]_23 ;
  wire [3:0]\reg_entries_0_reg[4]_24 ;
  wire \reg_entries_0_reg[4]_25 ;
  wire [1:0]\reg_entries_0_reg[4]_3 ;
  wire [1:0]\reg_entries_0_reg[4]_4 ;
  wire [3:0]\reg_entries_0_reg[4]_5 ;
  wire [3:0]\reg_entries_0_reg[4]_6 ;
  wire [3:0]\reg_entries_0_reg[4]_7 ;
  wire \reg_entries_0_reg[4]_8 ;
  wire [3:0]\reg_entries_0_reg[4]_9 ;
  wire [0:0]\reg_entries_0_reg[5] ;
  wire [3:0]\reg_entries_0_reg[5]_0 ;
  wire [3:0]\reg_entries_0_reg[5]_1 ;
  wire [2:0]\reg_entries_0_reg[5]_10 ;
  wire [2:0]\reg_entries_0_reg[5]_11 ;
  wire [2:0]\reg_entries_0_reg[5]_12 ;
  wire [2:0]\reg_entries_0_reg[5]_13 ;
  wire [2:0]\reg_entries_0_reg[5]_14 ;
  wire [2:0]\reg_entries_0_reg[5]_15 ;
  wire [3:0]\reg_entries_0_reg[5]_16 ;
  wire [3:0]\reg_entries_0_reg[5]_17 ;
  wire [3:0]\reg_entries_0_reg[5]_18 ;
  wire [3:0]\reg_entries_0_reg[5]_19 ;
  wire [3:0]\reg_entries_0_reg[5]_2 ;
  wire [3:0]\reg_entries_0_reg[5]_20 ;
  wire [3:0]\reg_entries_0_reg[5]_21 ;
  wire [3:0]\reg_entries_0_reg[5]_22 ;
  wire [3:0]\reg_entries_0_reg[5]_23 ;
  wire [3:0]\reg_entries_0_reg[5]_24 ;
  wire [3:0]\reg_entries_0_reg[5]_25 ;
  wire [0:0]\reg_entries_0_reg[5]_26 ;
  wire [3:0]\reg_entries_0_reg[5]_27 ;
  wire [3:0]\reg_entries_0_reg[5]_28 ;
  wire [0:0]\reg_entries_0_reg[5]_29 ;
  wire [3:0]\reg_entries_0_reg[5]_3 ;
  wire [3:0]\reg_entries_0_reg[5]_30 ;
  wire [3:0]\reg_entries_0_reg[5]_31 ;
  wire [0:0]\reg_entries_0_reg[5]_32 ;
  wire [3:0]\reg_entries_0_reg[5]_33 ;
  wire [3:0]\reg_entries_0_reg[5]_34 ;
  wire [0:0]\reg_entries_0_reg[5]_35 ;
  wire [3:0]\reg_entries_0_reg[5]_36 ;
  wire [3:0]\reg_entries_0_reg[5]_37 ;
  wire [0:0]\reg_entries_0_reg[5]_38 ;
  wire [3:0]\reg_entries_0_reg[5]_39 ;
  wire [3:0]\reg_entries_0_reg[5]_4 ;
  wire [3:0]\reg_entries_0_reg[5]_40 ;
  wire [0:0]\reg_entries_0_reg[5]_41 ;
  wire [3:0]\reg_entries_0_reg[5]_42 ;
  wire [3:0]\reg_entries_0_reg[5]_43 ;
  wire [0:0]\reg_entries_0_reg[5]_44 ;
  wire [3:0]\reg_entries_0_reg[5]_45 ;
  wire [3:0]\reg_entries_0_reg[5]_46 ;
  wire [0:0]\reg_entries_0_reg[5]_47 ;
  wire [3:0]\reg_entries_0_reg[5]_5 ;
  wire [3:0]\reg_entries_0_reg[5]_6 ;
  wire [3:0]\reg_entries_0_reg[5]_7 ;
  wire [2:0]\reg_entries_0_reg[5]_8 ;
  wire [2:0]\reg_entries_0_reg[5]_9 ;
  wire [2:0]\reg_entries_0_reg[6] ;
  wire [2:0]\reg_entries_0_reg[6]_0 ;
  wire \reg_entries_0_reg[6]_1 ;
  wire [2:0]\reg_entries_0_reg[6]_10 ;
  wire [2:0]\reg_entries_0_reg[6]_11 ;
  wire [2:0]\reg_entries_0_reg[6]_12 ;
  wire [2:0]\reg_entries_0_reg[6]_13 ;
  wire [0:0]\reg_entries_0_reg[6]_14 ;
  wire [1:0]\reg_entries_0_reg[6]_15 ;
  wire [1:0]\reg_entries_0_reg[6]_16 ;
  wire [1:0]\reg_entries_0_reg[6]_17 ;
  wire [3:0]\reg_entries_0_reg[6]_18 ;
  wire [3:0]\reg_entries_0_reg[6]_19 ;
  wire \reg_entries_0_reg[6]_2 ;
  wire [3:0]\reg_entries_0_reg[6]_20 ;
  wire [3:0]\reg_entries_0_reg[6]_21 ;
  wire [3:0]\reg_entries_0_reg[6]_22 ;
  wire [3:0]\reg_entries_0_reg[6]_23 ;
  wire [3:0]\reg_entries_0_reg[6]_24 ;
  wire [3:0]\reg_entries_0_reg[6]_25 ;
  wire [3:0]\reg_entries_0_reg[6]_26 ;
  wire [2:0]\reg_entries_0_reg[6]_27 ;
  wire [3:0]\reg_entries_0_reg[6]_28 ;
  wire [3:0]\reg_entries_0_reg[6]_29 ;
  wire \reg_entries_0_reg[6]_3 ;
  wire [3:0]\reg_entries_0_reg[6]_30 ;
  wire [3:0]\reg_entries_0_reg[6]_31 ;
  wire [3:0]\reg_entries_0_reg[6]_32 ;
  wire [3:0]\reg_entries_0_reg[6]_33 ;
  wire [3:0]\reg_entries_0_reg[6]_34 ;
  wire [3:0]\reg_entries_0_reg[6]_35 ;
  wire [3:0]\reg_entries_0_reg[6]_36 ;
  wire [3:0]\reg_entries_0_reg[6]_37 ;
  wire [2:0]\reg_entries_0_reg[6]_38 ;
  wire [3:0]\reg_entries_0_reg[6]_39 ;
  wire \reg_entries_0_reg[6]_4 ;
  wire [2:0]\reg_entries_0_reg[6]_40 ;
  wire [2:0]\reg_entries_0_reg[6]_41 ;
  wire \reg_entries_0_reg[6]_42 ;
  wire [3:0]\reg_entries_0_reg[6]_43 ;
  wire [3:0]\reg_entries_0_reg[6]_44 ;
  wire \reg_entries_0_reg[6]_45 ;
  wire [3:0]\reg_entries_0_reg[6]_46 ;
  wire [3:0]\reg_entries_0_reg[6]_47 ;
  wire \reg_entries_0_reg[6]_48 ;
  wire [3:0]\reg_entries_0_reg[6]_49 ;
  wire [1:0]\reg_entries_0_reg[6]_5 ;
  wire [3:0]\reg_entries_0_reg[6]_50 ;
  wire [3:0]\reg_entries_0_reg[6]_51 ;
  wire [3:0]\reg_entries_0_reg[6]_52 ;
  wire \reg_entries_0_reg[6]_53 ;
  wire [3:0]\reg_entries_0_reg[6]_54 ;
  wire [3:0]\reg_entries_0_reg[6]_55 ;
  wire [3:0]\reg_entries_0_reg[6]_56 ;
  wire [3:0]\reg_entries_0_reg[6]_57 ;
  wire \reg_entries_0_reg[6]_6 ;
  wire \reg_entries_0_reg[6]_7 ;
  wire [2:0]\reg_entries_0_reg[6]_8 ;
  wire [2:0]\reg_entries_0_reg[6]_9 ;
  wire \reg_entries_1_reg[0] ;
  wire \reg_entries_1_reg[0]_0 ;
  wire \reg_entries_1_reg[0]_1 ;
  wire [2:0]\reg_entries_1_reg[0]_10 ;
  wire [2:0]\reg_entries_1_reg[0]_11 ;
  wire [2:0]\reg_entries_1_reg[0]_12 ;
  wire [2:0]\reg_entries_1_reg[0]_13 ;
  wire [2:0]\reg_entries_1_reg[0]_14 ;
  wire \reg_entries_1_reg[0]_15 ;
  wire \reg_entries_1_reg[0]_16 ;
  wire \reg_entries_1_reg[0]_17 ;
  wire \reg_entries_1_reg[0]_18 ;
  wire \reg_entries_1_reg[0]_19 ;
  wire \reg_entries_1_reg[0]_2 ;
  wire \reg_entries_1_reg[0]_20 ;
  wire \reg_entries_1_reg[0]_21 ;
  wire \reg_entries_1_reg[0]_22 ;
  wire \reg_entries_1_reg[0]_23 ;
  wire \reg_entries_1_reg[0]_24 ;
  wire \reg_entries_1_reg[0]_25 ;
  wire \reg_entries_1_reg[0]_26 ;
  wire \reg_entries_1_reg[0]_27 ;
  wire \reg_entries_1_reg[0]_28 ;
  wire \reg_entries_1_reg[0]_29 ;
  wire \reg_entries_1_reg[0]_3 ;
  wire \reg_entries_1_reg[0]_30 ;
  wire \reg_entries_1_reg[0]_31 ;
  wire [0:0]\reg_entries_1_reg[0]_32 ;
  wire [0:0]\reg_entries_1_reg[0]_33 ;
  wire [0:0]\reg_entries_1_reg[0]_34 ;
  wire [0:0]\reg_entries_1_reg[0]_35 ;
  wire [0:0]\reg_entries_1_reg[0]_36 ;
  wire [0:0]\reg_entries_1_reg[0]_37 ;
  wire [0:0]\reg_entries_1_reg[0]_38 ;
  wire [0:0]\reg_entries_1_reg[0]_39 ;
  wire \reg_entries_1_reg[0]_4 ;
  wire [0:0]\reg_entries_1_reg[0]_40 ;
  wire [0:0]\reg_entries_1_reg[0]_41 ;
  wire [0:0]\reg_entries_1_reg[0]_42 ;
  wire [0:0]\reg_entries_1_reg[0]_43 ;
  wire [0:0]\reg_entries_1_reg[0]_44 ;
  wire [0:0]\reg_entries_1_reg[0]_45 ;
  wire [0:0]\reg_entries_1_reg[0]_46 ;
  wire [0:0]\reg_entries_1_reg[0]_47 ;
  wire \reg_entries_1_reg[0]_5 ;
  wire \reg_entries_1_reg[0]_6 ;
  wire \reg_entries_1_reg[0]_7 ;
  wire [2:0]\reg_entries_1_reg[0]_8 ;
  wire \reg_entries_1_reg[0]_9 ;
  wire [0:0]\reg_entries_1_reg[12] ;
  wire [2:0]\reg_entries_2_reg[12] ;
  wire [0:0]\reg_entries_3_reg[11] ;
  wire [2:0]\reg_entries_3_reg[12] ;
  wire [9:0]\reg_entries_4_reg[61] ;
  wire \reg_entries_4_reg[61]_0 ;
  wire \reg_mbadaddr_reg[12] ;
  wire \reg_mcause_reg[0] ;
  wire \reg_mepc_reg[12] ;
  wire [0:0]\reg_mie_reg[7] ;
  wire reg_mip_seip_reg;
  wire reg_mip_seip_reg_0;
  wire \reg_misa_reg[0] ;
  wire [1:0]\reg_misa_reg[12] ;
  wire \reg_misa_reg[12]_0 ;
  wire reg_mstatus_mie;
  wire reg_mstatus_mie_reg;
  wire reg_mstatus_mie_reg_0;
  wire reg_mstatus_mpie_reg;
  wire reg_mstatus_mpie_reg_0;
  wire \reg_mstatus_mpp_reg[0] ;
  wire \reg_mstatus_mpp_reg[1] ;
  wire \reg_mstatus_prv_reg[1] ;
  wire \reg_mstatus_prv_reg[1]_0 ;
  wire \reg_mstatus_prv_reg[1]_1 ;
  wire \reg_mstatus_prv_reg[1]_2 ;
  wire reg_mstatus_spie_reg;
  wire reg_mstatus_tvm_reg;
  wire \reg_mtvec_reg[10] ;
  wire \reg_mtvec_reg[11] ;
  wire \reg_mtvec_reg[12] ;
  wire \reg_mtvec_reg[13] ;
  wire \reg_mtvec_reg[14] ;
  wire \reg_mtvec_reg[15] ;
  wire \reg_mtvec_reg[16] ;
  wire \reg_mtvec_reg[17] ;
  wire \reg_mtvec_reg[18] ;
  wire \reg_mtvec_reg[19] ;
  wire \reg_mtvec_reg[20] ;
  wire \reg_mtvec_reg[20]_0 ;
  wire \reg_mtvec_reg[21] ;
  wire \reg_mtvec_reg[21]_0 ;
  wire \reg_mtvec_reg[22] ;
  wire \reg_mtvec_reg[22]_0 ;
  wire \reg_mtvec_reg[23] ;
  wire \reg_mtvec_reg[24] ;
  wire \reg_mtvec_reg[25] ;
  wire \reg_mtvec_reg[26] ;
  wire \reg_mtvec_reg[27] ;
  wire \reg_mtvec_reg[28] ;
  wire [28:0]\reg_mtvec_reg[29] ;
  wire [29:0]\reg_mtvec_reg[29]_0 ;
  wire [27:0]\reg_mtvec_reg[29]_1 ;
  wire [29:0]\reg_mtvec_reg[29]_2 ;
  wire [29:0]\reg_mtvec_reg[29]_3 ;
  wire [27:0]\reg_mtvec_reg[29]_4 ;
  wire [28:0]\reg_mtvec_reg[29]_5 ;
  wire [28:0]\reg_mtvec_reg[29]_6 ;
  wire \reg_mtvec_reg[29]_7 ;
  wire \reg_mtvec_reg[30] ;
  wire \reg_mtvec_reg[31] ;
  wire \reg_mtvec_reg[4] ;
  wire \reg_mtvec_reg[8] ;
  wire \reg_pmp_0_addr_reg[13] ;
  wire \reg_pmp_0_addr_reg[17] ;
  wire \reg_pmp_0_addr_reg[19] ;
  wire \reg_pmp_0_addr_reg[23] ;
  wire [0:0]\reg_pmp_0_addr_reg[28] ;
  wire [0:0]\reg_pmp_0_addr_reg[28]_0 ;
  wire \reg_pmp_0_addr_reg[29] ;
  wire [0:0]\reg_pmp_0_addr_reg[29]_0 ;
  wire \reg_pmp_1_addr_reg[13] ;
  wire \reg_pmp_1_addr_reg[17] ;
  wire \reg_pmp_1_addr_reg[19] ;
  wire [0:0]\reg_pmp_1_addr_reg[28] ;
  wire [0:0]\reg_pmp_1_addr_reg[28]_0 ;
  wire \reg_pmp_1_addr_reg[29] ;
  wire [0:0]\reg_pmp_1_addr_reg[29]_0 ;
  wire \reg_pmp_1_cfg_a_reg[0] ;
  wire reg_pmp_1_cfg_w_reg;
  wire \reg_pmp_2_addr_reg[0] ;
  wire \reg_pmp_2_addr_reg[13] ;
  wire \reg_pmp_2_addr_reg[17] ;
  wire \reg_pmp_2_addr_reg[19] ;
  wire [0:0]\reg_pmp_2_addr_reg[28] ;
  wire [0:0]\reg_pmp_2_addr_reg[28]_0 ;
  wire \reg_pmp_2_addr_reg[29] ;
  wire \reg_pmp_2_addr_reg[29]_0 ;
  wire [0:0]\reg_pmp_2_addr_reg[29]_1 ;
  wire \reg_pmp_2_cfg_a_reg[0] ;
  wire \reg_pmp_3_addr_reg[13] ;
  wire \reg_pmp_3_addr_reg[17] ;
  wire \reg_pmp_3_addr_reg[18] ;
  wire \reg_pmp_3_addr_reg[19] ;
  wire \reg_pmp_3_addr_reg[23] ;
  wire [0:0]\reg_pmp_3_addr_reg[28] ;
  wire [0:0]\reg_pmp_3_addr_reg[28]_0 ;
  wire \reg_pmp_3_addr_reg[29] ;
  wire [0:0]\reg_pmp_3_addr_reg[29]_0 ;
  wire \reg_pmp_3_addr_reg[29]_1 ;
  wire \reg_pmp_4_addr_reg[0] ;
  wire \reg_pmp_4_addr_reg[13] ;
  wire \reg_pmp_4_addr_reg[14] ;
  wire \reg_pmp_4_addr_reg[17] ;
  wire \reg_pmp_4_addr_reg[19] ;
  wire [0:0]\reg_pmp_4_addr_reg[28] ;
  wire [0:0]\reg_pmp_4_addr_reg[28]_0 ;
  wire \reg_pmp_4_addr_reg[29] ;
  wire [0:0]\reg_pmp_4_addr_reg[29]_0 ;
  wire [0:0]\reg_pmp_4_cfg_a_reg[1] ;
  wire \reg_pmp_5_addr_reg[13] ;
  wire \reg_pmp_5_addr_reg[17] ;
  wire \reg_pmp_5_addr_reg[19] ;
  wire \reg_pmp_5_addr_reg[20] ;
  wire [0:0]\reg_pmp_5_addr_reg[28] ;
  wire [0:0]\reg_pmp_5_addr_reg[28]_0 ;
  wire \reg_pmp_5_addr_reg[29] ;
  wire [0:0]\reg_pmp_5_addr_reg[29]_0 ;
  wire [0:0]\reg_pmp_5_cfg_a_reg[1] ;
  wire \reg_pmp_5_cfg_a_reg[1]_0 ;
  wire \reg_pmp_6_addr_reg[13] ;
  wire \reg_pmp_6_addr_reg[17] ;
  wire \reg_pmp_6_addr_reg[19] ;
  wire [0:0]\reg_pmp_6_addr_reg[28] ;
  wire [0:0]\reg_pmp_6_addr_reg[28]_0 ;
  wire \reg_pmp_6_addr_reg[29] ;
  wire [0:0]\reg_pmp_6_addr_reg[29]_0 ;
  wire \reg_pmp_7_addr_reg[13] ;
  wire \reg_pmp_7_addr_reg[17] ;
  wire \reg_pmp_7_addr_reg[17]_0 ;
  wire \reg_pmp_7_addr_reg[19] ;
  wire \reg_pmp_7_addr_reg[23] ;
  wire [0:0]\reg_pmp_7_addr_reg[28] ;
  wire [0:0]\reg_pmp_7_addr_reg[28]_0 ;
  wire \reg_pmp_7_addr_reg[29] ;
  wire \reg_pmp_7_addr_reg[29]_0 ;
  wire [0:0]\reg_pmp_7_addr_reg[29]_1 ;
  wire \reg_pmp_7_addr_reg[29]_2 ;
  wire \reg_pmp_7_cfg_a_reg[0] ;
  wire \reg_sbadaddr_reg[0] ;
  wire [2:0]\reg_sbadaddr_reg[30] ;
  wire [2:0]\reg_sbadaddr_reg[30]_0 ;
  wire [2:0]\reg_sbadaddr_reg[30]_1 ;
  wire [1:0]\reg_sbadaddr_reg[30]_2 ;
  wire \reg_sbadaddr_reg[30]_3 ;
  wire [2:0]\reg_sbadaddr_reg[30]_4 ;
  wire [1:0]\reg_sbadaddr_reg[30]_5 ;
  wire [2:0]\reg_sbadaddr_reg[30]_6 ;
  wire [1:0]\reg_sbadaddr_reg[30]_7 ;
  wire [1:0]\reg_sbadaddr_reg[30]_8 ;
  wire [1:0]\reg_sbadaddr_reg[30]_9 ;
  wire [0:0]\reg_sbadaddr_reg[39] ;
  wire [0:0]\reg_sbadaddr_reg[39]_0 ;
  wire [3:0]\reg_sbadaddr_reg[39]_1 ;
  wire [3:0]\reg_sbadaddr_reg[39]_2 ;
  wire \reg_scause_reg[0] ;
  wire \reg_scause_reg[0]_0 ;
  wire \reg_scause_reg[1] ;
  wire \reg_scause_reg[1]_0 ;
  wire [0:0]\reg_scause_reg[2] ;
  wire \reg_scause_reg[3] ;
  wire \reg_sepc_reg[12] ;
  wire \reg_sepc_reg[26] ;
  wire reg_singleStepped;
  wire \reg_sptbr_ppn[19]_i_4_n_0 ;
  wire \reg_sptbr_ppn_reg[0] ;
  wire \reg_sscratch_reg[0] ;
  wire [4:0]\reg_sscratch_reg[45] ;
  wire \reg_sscratch_reg[45]_0 ;
  wire [2:0]\reg_sscratch_reg[59] ;
  wire [23:0]\reg_sscratch_reg[62] ;
  wire \reg_stvec_reg[32] ;
  wire \reg_stvec_reg[33] ;
  wire \reg_stvec_reg[34] ;
  wire \reg_stvec_reg[35] ;
  wire \reg_stvec_reg[36] ;
  wire \reg_stvec_reg[37] ;
  wire \reg_stvec_reg[38] ;
  wire reg_wfi_reg;
  wire [3:0]\remainder_reg[103] ;
  wire [0:0]\remainder_reg[103]_0 ;
  wire [2:0]\remainder_reg[103]_1 ;
  wire [3:0]\remainder_reg[103]_2 ;
  wire [3:0]\remainder_reg[107] ;
  wire [3:0]\remainder_reg[107]_0 ;
  wire [3:0]\remainder_reg[107]_1 ;
  wire [3:0]\remainder_reg[111] ;
  wire [3:0]\remainder_reg[111]_0 ;
  wire [3:0]\remainder_reg[111]_1 ;
  wire [3:0]\remainder_reg[115] ;
  wire [0:0]\remainder_reg[115]_0 ;
  wire [2:0]\remainder_reg[115]_1 ;
  wire [3:0]\remainder_reg[115]_2 ;
  wire [3:0]\remainder_reg[119] ;
  wire [3:0]\remainder_reg[119]_0 ;
  wire [3:0]\remainder_reg[123] ;
  wire [3:0]\remainder_reg[123]_0 ;
  wire [0:0]\remainder_reg[127] ;
  wire [3:0]\remainder_reg[127]_0 ;
  wire [3:0]\remainder_reg[127]_1 ;
  wire [3:0]\remainder_reg[127]_2 ;
  wire [1:0]\remainder_reg[127]_3 ;
  wire [3:0]\remainder_reg[127]_4 ;
  wire [3:0]\remainder_reg[127]_5 ;
  wire [0:0]\remainder_reg[127]_6 ;
  wire [3:0]\remainder_reg[127]_7 ;
  wire [0:0]\remainder_reg[128] ;
  wire \remainder_reg[129] ;
  wire \remainder_reg[129]_0 ;
  wire [2:0]\remainder_reg[129]_1 ;
  wire \remainder_reg[31] ;
  wire \remainder_reg[33] ;
  wire \remainder_reg[33]_0 ;
  wire \remainder_reg[34] ;
  wire \remainder_reg[34]_0 ;
  wire \remainder_reg[35] ;
  wire \remainder_reg[35]_0 ;
  wire \remainder_reg[36] ;
  wire \remainder_reg[36]_0 ;
  wire \remainder_reg[37] ;
  wire \remainder_reg[37]_0 ;
  wire \remainder_reg[38] ;
  wire \remainder_reg[38]_0 ;
  wire \remainder_reg[39] ;
  wire \remainder_reg[41] ;
  wire \remainder_reg[42] ;
  wire \remainder_reg[43] ;
  wire \remainder_reg[44] ;
  wire \remainder_reg[46] ;
  wire \remainder_reg[47] ;
  wire \remainder_reg[49] ;
  wire \remainder_reg[50] ;
  wire \remainder_reg[51] ;
  wire \remainder_reg[52] ;
  wire \remainder_reg[54] ;
  wire \remainder_reg[55] ;
  wire \remainder_reg[57] ;
  wire \remainder_reg[58] ;
  wire \remainder_reg[59] ;
  wire \remainder_reg[60] ;
  wire \remainder_reg[61] ;
  wire \remainder_reg[62] ;
  wire [24:0]\remainder_reg[62]_0 ;
  wire \remainder_reg[63] ;
  wire [2:0]\remainder_reg[64] ;
  wire [3:0]\remainder_reg[64]_0 ;
  wire [3:0]\remainder_reg[64]_1 ;
  wire [2:0]\remainder_reg[64]_2 ;
  wire [2:0]\remainder_reg[64]_3 ;
  wire [3:0]\remainder_reg[64]_4 ;
  wire [3:0]\remainder_reg[64]_5 ;
  wire [3:0]\remainder_reg[64]_6 ;
  wire [0:0]\remainder_reg[64]_7 ;
  wire [3:0]\remainder_reg[64]_8 ;
  wire [0:0]\remainder_reg[64]_9 ;
  wire [64:0]\remainder_reg[65] ;
  wire [3:0]\remainder_reg[71] ;
  wire [3:0]\remainder_reg[75] ;
  wire [3:0]\remainder_reg[79] ;
  wire [3:0]\remainder_reg[83] ;
  wire [3:0]\remainder_reg[87] ;
  wire [3:0]\remainder_reg[91] ;
  wire [3:0]\remainder_reg[91]_0 ;
  wire [3:0]\remainder_reg[95] ;
  wire [3:0]\remainder_reg[95]_0 ;
  wire [3:0]\remainder_reg[99] ;
  wire [3:0]\remainder_reg[99]_0 ;
  wire req_dw_reg;
  wire \req_tag_reg[0] ;
  wire \req_tag_reg[0]_0 ;
  wire \req_tag_reg[1] ;
  wire \req_tag_reg[1]_0 ;
  wire \req_tag_reg[1]_1 ;
  wire \req_tag_reg[1]_2 ;
  wire \req_tag_reg[1]_3 ;
  wire \req_tag_reg[1]_4 ;
  wire \req_tag_reg[4] ;
  wire resHi_reg;
  wire resp_valid_0_reg;
  wire resp_valid_1_reg;
  wire \s1_pc[10]_i_4_n_0 ;
  wire \s1_pc[11]_i_4_n_0 ;
  wire \s1_pc[12]_i_5_n_0 ;
  wire \s1_pc[13]_i_4_n_0 ;
  wire \s1_pc[14]_i_4_n_0 ;
  wire \s1_pc[15]_i_4_n_0 ;
  wire \s1_pc[16]_i_5_n_0 ;
  wire \s1_pc[17]_i_4_n_0 ;
  wire \s1_pc[18]_i_4_n_0 ;
  wire \s1_pc[19]_i_4_n_0 ;
  wire \s1_pc[1]_i_3_n_0 ;
  wire \s1_pc[20]_i_5_n_0 ;
  wire \s1_pc[21]_i_4_n_0 ;
  wire \s1_pc[22]_i_4_n_0 ;
  wire \s1_pc[23]_i_4_n_0 ;
  wire \s1_pc[24]_i_5_n_0 ;
  wire \s1_pc[25]_i_4_n_0 ;
  wire \s1_pc[26]_i_4_n_0 ;
  wire \s1_pc[27]_i_4_n_0 ;
  wire \s1_pc[28]_i_5_n_0 ;
  wire \s1_pc[29]_i_4_n_0 ;
  wire \s1_pc[2]_i_4_n_0 ;
  wire \s1_pc[30]_i_4_n_0 ;
  wire \s1_pc[31]_i_4_n_0 ;
  wire \s1_pc[32]_i_4_n_0 ;
  wire \s1_pc[33]_i_3_n_0 ;
  wire \s1_pc[34]_i_3_n_0 ;
  wire \s1_pc[35]_i_3_n_0 ;
  wire \s1_pc[36]_i_4_n_0 ;
  wire \s1_pc[37]_i_3_n_0 ;
  wire \s1_pc[38]_i_3_n_0 ;
  wire \s1_pc[39]_i_4_n_0 ;
  wire \s1_pc[3]_i_4_n_0 ;
  wire \s1_pc[3]_i_7_n_0 ;
  wire \s1_pc[4]_i_4_n_0 ;
  wire \s1_pc[5]_i_3_n_0 ;
  wire \s1_pc[6]_i_4_n_0 ;
  wire \s1_pc[7]_i_4_n_0 ;
  wire \s1_pc[8]_i_5_n_0 ;
  wire \s1_pc[9]_i_4_n_0 ;
  wire [0:0]\s1_pc_reg[1] ;
  wire \s1_pc_reg[26] ;
  wire \s1_pc_reg[31] ;
  wire [37:0]\s1_pc_reg[39]_0 ;
  wire [3:0]\s1_pc_reg[39]_1 ;
  wire [3:0]\s1_pc_reg[39]_2 ;
  wire [3:0]\s1_pc_reg[39]_3 ;
  wire [3:0]\s1_pc_reg[39]_4 ;
  wire [0:0]\s1_pc_reg[39]_5 ;
  wire [11:0]\s1_pc_reg[39]_6 ;
  wire [0:0]\s1_pc_reg[4] ;
  wire [0:0]\s1_pc_reg[4]_0 ;
  wire \s1_pc_reg[5] ;
  wire \s1_req_addr_reg[2] ;
  wire \s1_req_addr_reg[2]_0 ;
  wire \s1_req_addr_reg[2]_1 ;
  wire \s1_req_addr_reg[2]_2 ;
  wire [10:0]\s1_req_addr_reg[31] ;
  wire [18:0]\s1_req_addr_reg[39] ;
  wire [3:0]\s1_req_addr_reg[39]_0 ;
  wire [3:0]\s1_req_addr_reg[39]_1 ;
  wire [3:0]\s1_req_addr_reg[39]_2 ;
  wire [3:0]\s1_req_addr_reg[39]_3 ;
  wire [0:0]\s1_req_addr_reg[39]_4 ;
  wire [0:0]\s1_req_addr_reg[3] ;
  wire [4:0]\s1_req_cmd_reg[4] ;
  wire s1_req_phys_reg;
  wire s1_req_phys_reg_0;
  wire \s1_req_typ_reg[0] ;
  wire \s1_req_typ_reg[0]_0 ;
  wire \s1_req_typ_reg[0]_1 ;
  wire \s1_req_typ_reg[0]_2 ;
  wire \s1_req_typ_reg[0]_3 ;
  wire \s1_req_typ_reg[1] ;
  wire s1_valid_reg;
  wire [0:0]\s2_pc_reg[1] ;
  wire s2_replay;
  wire [1:0]\s2_req_addr_reg[31] ;
  wire \s2_req_cmd_reg[1] ;
  wire \s2_req_tag_reg[5] ;
  wire \s2_req_tag_reg[5]_0 ;
  wire [4:0]\s2_req_tag_reg[6] ;
  wire \s2_req_tag_reg[6]_0 ;
  wire [19:0]\s2_req_typ_reg[0] ;
  wire s2_tlb_resp_cacheable_reg;
  wire s2_valid_reg;
  wire [0:0]shamt;
  wire \state_reg[0] ;
  wire \state_reg[0]_0 ;
  wire \state_reg[0]_1 ;
  wire \state_reg[0]_2 ;
  wire \state_reg[1] ;
  wire \state_reg[1]_0 ;
  wire \state_reg[1]_1 ;
  wire \state_reg[2] ;
  wire sys_reset_reg;
  wire sys_reset_reg_0;
  wire sys_reset_reg_1;
  wire sys_reset_reg_2;
  wire target_reset;
  wire tile_auto_int_sync_xing_sinklzy_in_0_sync_0;
  wire tile_auto_int_sync_xing_sinklzy_in_0_sync_1;
  wire tile_auto_int_sync_xing_sinklzy_in_1_sync_0;
  wire tile_auto_int_sync_xing_sinklzy_in_2_sync_0;
  wire tlb_io_req_bits_sfence_bits_rs2;
  wire trig_jalr_count;
  wire \trig_jalr_count[4]_i_3_n_0 ;
  wire \trig_jalr_count[4]_i_4_n_0 ;
  wire \trig_jalr_count_reg[0]_0 ;
  wire [3:0]\trig_jalr_count_reg[0]_1 ;
  wire [3:0]\trig_jalr_count_reg[0]_2 ;
  wire [3:0]\trig_jalr_count_reg[0]_3 ;
  wire [3:0]\trig_jalr_count_reg[0]_4 ;
  wire [3:0]\trig_jalr_count_reg[0]_5 ;
  wire [0:0]\trig_jalr_count_reg[0]_6 ;
  wire [4:0]trig_jalr_count_reg__0;
  wire \trig_mem_data[120]_i_1_n_0 ;
  wire \trig_mem_data[125]_i_1_n_0 ;
  wire \trig_mem_data[126]_i_1_n_0 ;
  wire \trig_mem_data[127]_i_10_n_0 ;
  wire \trig_mem_data[127]_i_11_n_0 ;
  wire \trig_mem_data[127]_i_12_n_0 ;
  wire \trig_mem_data[127]_i_13_n_0 ;
  wire \trig_mem_data[127]_i_14_n_0 ;
  wire \trig_mem_data[127]_i_15_n_0 ;
  wire \trig_mem_data[127]_i_2_n_0 ;
  wire \trig_mem_data[127]_i_3_n_0 ;
  wire \trig_mem_data[127]_i_4_n_0 ;
  wire \trig_mem_data[127]_i_5_n_0 ;
  wire \trig_mem_data[127]_i_6_n_0 ;
  wire \trig_mem_data[127]_i_7_n_0 ;
  wire \trig_mem_data[127]_i_8_n_0 ;
  wire \trig_mem_data[127]_i_9_n_0 ;
  wire [1:0]\trig_mem_data_reg[126]_0 ;
  wire [0:0]\trig_mem_data_reg[127]_0 ;
  wire [0:0]\trig_mem_data_reg[63]_0 ;
  wire \trig_mem_data_reg_n_0_[0] ;
  wire trig_pc;
  wire \trig_pc[0]_i_1_n_0 ;
  wire \trig_pc_reg[0]_0 ;
  wire \trig_pc_reg[0]_1 ;
  wire [3:0]\trig_pc_reg[0]_2 ;
  wire [3:0]\trig_pc_reg[0]_3 ;
  wire [3:0]\trig_pc_reg[0]_4 ;
  wire [3:0]\trig_pc_reg[0]_5 ;
  wire [3:0]\trig_pc_reg[0]_6 ;
  wire [0:0]\trig_pc_reg[0]_7 ;
  wire [63:0]\trig_pc_reg[63]_0 ;
  wire [0:0]\trig_pc_reg[63]_1 ;
  wire trig_pc_valid_reg_0;
  wire trig_pc_valid_reg_1;
  wire trig_pc_valid_reg_2;
  wire [0:0]trig_state;
  wire \trig_state[0]_i_1_n_0 ;
  wire \trig_state[0]_i_2_n_0 ;
  wire \trig_state[0]_i_4_n_0 ;
  wire \trig_state[1]_i_1_n_0 ;
  wire \trig_state[1]_i_2_n_0 ;
  wire \trig_state[1]_i_4_n_0 ;
  wire \trig_state_reg[0]_0 ;
  wire \trig_state_reg[0]_1 ;
  wire \trig_state_reg[1]_0 ;
  wire \trig_state_reg[1]_1 ;
  wire \trig_state_reg[1]_2 ;
  wire [3:0]\trig_state_reg[1]_3 ;
  wire [3:0]\trig_state_reg[1]_4 ;
  wire [3:0]\trig_state_reg[1]_5 ;
  wire [3:0]\trig_state_reg[1]_6 ;
  wire [3:0]\trig_state_reg[1]_7 ;
  wire [0:0]\trig_state_reg[1]_8 ;
  wire \valid_reg[0] ;
  wire \valid_reg[0]_0 ;
  wire \valid_reg[1] ;
  wire \valid_reg[1]_0 ;
  wire \valid_reg[2] ;
  wire \valid_reg[3] ;
  wire [0:0]\valid_reg[3]_0 ;
  wire [0:0]\valid_reg[3]_1 ;
  wire [0:0]\valid_reg[3]_2 ;
  wire \valid_reg[3]_3 ;
  wire [0:0]\valid_reg[3]_4 ;
  wire \valid_reg[4] ;
  wire \wb_ctrl_csr_reg[0]_0 ;
  wire [0:0]\wb_ctrl_csr_reg[0]_1 ;
  wire \wb_ctrl_csr_reg[0]_10 ;
  wire [0:0]\wb_ctrl_csr_reg[0]_2 ;
  wire [39:0]\wb_ctrl_csr_reg[0]_3 ;
  wire [0:0]\wb_ctrl_csr_reg[0]_4 ;
  wire [4:0]\wb_ctrl_csr_reg[0]_5 ;
  wire [0:0]\wb_ctrl_csr_reg[0]_6 ;
  wire [0:0]\wb_ctrl_csr_reg[0]_7 ;
  wire [5:0]\wb_ctrl_csr_reg[0]_8 ;
  wire [0:0]\wb_ctrl_csr_reg[0]_9 ;
  wire \wb_ctrl_csr_reg[2]_0 ;
  wire wb_ctrl_div;
  wire wb_ctrl_fence_i;
  wire wb_ctrl_fence_i_reg_0;
  wire wb_ctrl_mem;
  wire wb_ctrl_mem_reg_0;
  wire wb_ctrl_wxd;
  wire [63:0]wb_reg_cause;
  wire \wb_reg_cause[63]_i_1_n_0 ;
  wire \wb_reg_cause_reg[0]_0 ;
  wire [3:0]\wb_reg_cause_reg[0]_1 ;
  wire [3:0]\wb_reg_cause_reg[0]_10 ;
  wire [3:0]\wb_reg_cause_reg[0]_11 ;
  wire [3:0]\wb_reg_cause_reg[0]_12 ;
  wire [2:0]\wb_reg_cause_reg[0]_13 ;
  wire [2:0]\wb_reg_cause_reg[0]_14 ;
  wire [3:0]\wb_reg_cause_reg[0]_2 ;
  wire [3:0]\wb_reg_cause_reg[0]_3 ;
  wire [0:0]\wb_reg_cause_reg[0]_4 ;
  wire [3:0]\wb_reg_cause_reg[0]_5 ;
  wire [3:0]\wb_reg_cause_reg[0]_6 ;
  wire [3:0]\wb_reg_cause_reg[0]_7 ;
  wire [3:0]\wb_reg_cause_reg[0]_8 ;
  wire [3:0]\wb_reg_cause_reg[0]_9 ;
  wire \wb_reg_cause_reg[2]_0 ;
  wire [1:0]\wb_reg_cause_reg[3]_0 ;
  wire \wb_reg_cause_reg[63]_0 ;
  wire [0:0]\wb_reg_cause_reg[63]_1 ;
  wire [0:0]\wb_reg_cause_reg[63]_2 ;
  wire [0:0]\wb_reg_cause_reg[63]_3 ;
  wire [0:0]\wb_reg_cause_reg[63]_4 ;
  wire [0:0]\wb_reg_cause_reg[63]_5 ;
  wire [0:0]\wb_reg_cause_reg[63]_6 ;
  wire wb_reg_flush_pipe;
  wire wb_reg_flush_pipe0;
  wire \wb_reg_inst_reg[21]_0 ;
  wire \wb_reg_inst_reg[21]_1 ;
  wire \wb_reg_inst_reg[21]_2 ;
  wire \wb_reg_inst_reg[21]_3 ;
  wire \wb_reg_inst_reg[21]_4 ;
  wire \wb_reg_inst_reg[21]_5 ;
  wire \wb_reg_inst_reg[22]_0 ;
  wire \wb_reg_inst_reg[22]_1 ;
  wire \wb_reg_inst_reg[26]_0 ;
  wire \wb_reg_inst_reg[29]_0 ;
  wire \wb_reg_inst_reg[29]_1 ;
  wire \wb_reg_inst_reg[30]_0 ;
  wire \wb_reg_inst_reg[30]_1 ;
  wire [24:0]\wb_reg_inst_reg[31]_0 ;
  wire \wb_reg_inst_reg[7]_0 ;
  wire \wb_reg_inst_reg[7]_1 ;
  wire \wb_reg_inst_reg[9]_0 ;
  wire \wb_reg_inst_reg[9]_1 ;
  wire \wb_reg_inst_reg[9]_2 ;
  wire \wb_reg_inst_reg[9]_3 ;
  wire [3:0]\wb_reg_pc_reg[34]_0 ;
  wire [32:0]\wb_reg_pc_reg[39]_0 ;
  wire [38:0]\wb_reg_pc_reg[39]_1 ;
  wire [38:0]\wb_reg_pc_reg[39]_2 ;
  wire [38:0]\wb_reg_pc_reg[39]_3 ;
  wire wb_reg_replay;
  wire wb_reg_replay0;
  wire wb_reg_replay_reg_0;
  wire wb_reg_replay_reg_1;
  wire wb_reg_replay_reg_2;
  wire wb_reg_sfence;
  wire wb_reg_valid;
  wire wb_reg_valid_reg_0;
  wire wb_reg_xcpt;
  wire wb_reg_xcpt0;
  wire wb_reg_xcpt_i_2_n_0;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r1_0_31_0_5
       (.ADDRA(ADDRA),
        .ADDRB(ADDRA),
        .ADDRC(ADDRA),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[1:0]),
        .DIB(_GEN_274[3:2]),
        .DIC(_GEN_274[5:4]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1416),
        .DOB(_T_1416_0[3:2]),
        .DOC(_T_1416_0[5:4]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* SOFT_HLUTNM = "soft_lutpair1783" *) 
  LUT3 #(
    .INIT(8'h01)) 
    _T_1396_reg_r1_0_31_0_5_i_44
       (.I0(\reg_sscratch_reg[59] [2]),
        .I1(\reg_sscratch_reg[59] [0]),
        .I2(\reg_sscratch_reg[59] [1]),
        .O(_T_1396_reg_r1_0_31_0_5_i_44_n_0));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r1_0_31_12_17
       (.ADDRA(ADDRA),
        .ADDRB(ADDRA),
        .ADDRC(ADDRA),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(\s2_req_typ_reg[0] [3:2]),
        .DIB(\s2_req_typ_reg[0] [5:4]),
        .DIC(\s2_req_typ_reg[0] [7:6]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1416_0[13:12]),
        .DOB(_T_1416_0[15:14]),
        .DOC(_T_1416_0[17:16]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r1_0_31_18_23
       (.ADDRA(ADDRA),
        .ADDRB(ADDRA),
        .ADDRC(ADDRA),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(\s2_req_typ_reg[0] [9:8]),
        .DIB(\s2_req_typ_reg[0] [11:10]),
        .DIC(\s2_req_typ_reg[0] [13:12]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1416_0[19:18]),
        .DOB(_T_1416_0[21:20]),
        .DOC(_T_1416_0[23:22]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r1_0_31_24_29
       (.ADDRA(ADDRA),
        .ADDRB(ADDRA),
        .ADDRC(ADDRA),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(\s2_req_typ_reg[0] [15:14]),
        .DIB(\s2_req_typ_reg[0] [17:16]),
        .DIC(\s2_req_typ_reg[0] [19:18]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1416_0[25:24]),
        .DOB(_T_1416_0[27:26]),
        .DOC(_T_1416_0[29:28]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r1_0_31_30_35
       (.ADDRA(ADDRA),
        .ADDRB(ADDRA),
        .ADDRC(ADDRA),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[11:10]),
        .DIB(_GEN_274[13:12]),
        .DIC(_GEN_274[15:14]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1416_0[31:30]),
        .DOB(_T_1416_0[33:32]),
        .DOC(_T_1416_0[35:34]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r1_0_31_36_41
       (.ADDRA(ADDRA),
        .ADDRB(ADDRA),
        .ADDRC(ADDRA),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[17:16]),
        .DIB(_GEN_274[19:18]),
        .DIC(_GEN_274[21:20]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1416_0[37:36]),
        .DOB(_T_1416_0[39:38]),
        .DOC(_T_1416_0[41:40]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r1_0_31_42_47
       (.ADDRA(ADDRA),
        .ADDRB(ADDRA),
        .ADDRC(ADDRA),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[23:22]),
        .DIB(_GEN_274[25:24]),
        .DIC(_GEN_274[27:26]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1416_0[43:42]),
        .DOB(_T_1416_0[45:44]),
        .DOC(_T_1416_0[47:46]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r1_0_31_48_53
       (.ADDRA(ADDRA),
        .ADDRB(ADDRA),
        .ADDRC(ADDRA),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[29:28]),
        .DIB(_GEN_274[31:30]),
        .DIC(_GEN_274[33:32]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1416_0[49:48]),
        .DOB(_T_1416_0[51:50]),
        .DOC(_T_1416_0[53:52]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r1_0_31_54_59
       (.ADDRA(ADDRA),
        .ADDRB(ADDRA),
        .ADDRC(ADDRA),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[35:34]),
        .DIB(_GEN_274[37:36]),
        .DIC(_GEN_274[39:38]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1416_0[55:54]),
        .DOB(_T_1416_0[57:56]),
        .DOC(_T_1416_0[59:58]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r1_0_31_60_63
       (.ADDRA(ADDRA),
        .ADDRB(ADDRA),
        .ADDRC(ADDRA),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[41:40]),
        .DIB(_GEN_274[43:42]),
        .DIC({\<const0> ,\<const0> }),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1416_0[61:60]),
        .DOB(_T_1416_0[63:62]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r1_0_31_6_11
       (.ADDRA(ADDRA),
        .ADDRB(ADDRA),
        .ADDRC(ADDRA),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[7:6]),
        .DIB(_GEN_274[9:8]),
        .DIC(\s2_req_typ_reg[0] [1:0]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1416_0[7:6]),
        .DOB(_T_1416_0[9:8]),
        .DOC(_T_1416_0[11:10]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r2_0_31_0_5
       (.ADDRA(nBufValid_reg_6),
        .ADDRB(nBufValid_reg_6),
        .ADDRC(nBufValid_reg_6),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[1:0]),
        .DIB(_GEN_274[3:2]),
        .DIC(_GEN_274[5:4]),
        .DID({\<const0> ,\<const0> }),
        .DOA({_T_1406_1,_T_1406[0]}),
        .DOB(_T_1406[2:1]),
        .DOC(_T_1406[4:3]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r2_0_31_12_17
       (.ADDRA(nBufValid_reg_6),
        .ADDRB(nBufValid_reg_6),
        .ADDRC(nBufValid_reg_6),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(\s2_req_typ_reg[0] [3:2]),
        .DIB(\s2_req_typ_reg[0] [5:4]),
        .DIC(\s2_req_typ_reg[0] [7:6]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1406[12:11]),
        .DOB(_T_1406[14:13]),
        .DOC(_T_1406[16:15]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r2_0_31_18_23
       (.ADDRA(nBufValid_reg_6),
        .ADDRB(nBufValid_reg_6),
        .ADDRC(nBufValid_reg_6),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(\s2_req_typ_reg[0] [9:8]),
        .DIB(\s2_req_typ_reg[0] [11:10]),
        .DIC(\s2_req_typ_reg[0] [13:12]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1406[18:17]),
        .DOB(_T_1406[20:19]),
        .DOC(_T_1406[22:21]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r2_0_31_24_29
       (.ADDRA(nBufValid_reg_6),
        .ADDRB(nBufValid_reg_6),
        .ADDRC(nBufValid_reg_6),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(\s2_req_typ_reg[0] [15:14]),
        .DIB(\s2_req_typ_reg[0] [17:16]),
        .DIC(\s2_req_typ_reg[0] [19:18]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1406[24:23]),
        .DOB(_T_1406[26:25]),
        .DOC(_T_1406[28:27]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r2_0_31_30_35
       (.ADDRA(nBufValid_reg_6),
        .ADDRB(nBufValid_reg_6),
        .ADDRC(nBufValid_reg_6),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[11:10]),
        .DIB(_GEN_274[13:12]),
        .DIC(_GEN_274[15:14]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1406[30:29]),
        .DOB(_T_1406[32:31]),
        .DOC(_T_1406[34:33]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r2_0_31_36_41
       (.ADDRA(nBufValid_reg_6),
        .ADDRB(nBufValid_reg_6),
        .ADDRC(nBufValid_reg_6),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[17:16]),
        .DIB(_GEN_274[19:18]),
        .DIC(_GEN_274[21:20]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1406[36:35]),
        .DOB(_T_1406[38:37]),
        .DOC(_T_1406[40:39]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r2_0_31_42_47
       (.ADDRA(nBufValid_reg_6),
        .ADDRB(nBufValid_reg_6),
        .ADDRC(nBufValid_reg_6),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[23:22]),
        .DIB(_GEN_274[25:24]),
        .DIC(_GEN_274[27:26]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1406[42:41]),
        .DOB(_T_1406[44:43]),
        .DOC(_T_1406[46:45]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r2_0_31_48_53
       (.ADDRA(nBufValid_reg_6),
        .ADDRB(nBufValid_reg_6),
        .ADDRC(nBufValid_reg_6),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[29:28]),
        .DIB(_GEN_274[31:30]),
        .DIC(_GEN_274[33:32]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1406[48:47]),
        .DOB(_T_1406[50:49]),
        .DOC(_T_1406[52:51]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r2_0_31_54_59
       (.ADDRA(nBufValid_reg_6),
        .ADDRB(nBufValid_reg_6),
        .ADDRC(nBufValid_reg_6),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[35:34]),
        .DIB(_GEN_274[37:36]),
        .DIC(_GEN_274[39:38]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1406[54:53]),
        .DOB(_T_1406[56:55]),
        .DOC(_T_1406[58:57]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r2_0_31_60_63
       (.ADDRA(nBufValid_reg_6),
        .ADDRB(nBufValid_reg_6),
        .ADDRC(nBufValid_reg_6),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[41:40]),
        .DIB(_GEN_274[43:42]),
        .DIC({\<const0> ,\<const0> }),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1406[60:59]),
        .DOB(_T_1406[62:61]),
        .WCLK(host_clk),
        .WE(p_31_in));
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)) 
    _T_1396_reg_r2_0_31_6_11
       (.ADDRA(nBufValid_reg_6),
        .ADDRB(nBufValid_reg_6),
        .ADDRC(nBufValid_reg_6),
        .ADDRD({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        .DIA(_GEN_274[7:6]),
        .DIB(_GEN_274[9:8]),
        .DIC(\s2_req_typ_reg[0] [1:0]),
        .DID({\<const0> ,\<const0> }),
        .DOA(_T_1406[6:5]),
        .DOB(_T_1406[8:7]),
        .DOC(_T_1406[10:9]),
        .WCLK(host_clk),
        .WE(p_31_in));
  FDRE #(
    .INIT(1'b0)) 
    _T_2373_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ex_ctrl_div_reg_0),
        .Q(_T_2373),
        .R(\<const0> ));
  (* SOFT_HLUTNM = "soft_lutpair1877" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \_T_2547[15]_i_3 
       (.I0(\reg_bp_0_control_tmatch_reg[1] [4]),
        .I1(\_T_2547[31]_i_6_n_0 ),
        .I2(\reg_bp_0_control_tmatch_reg[1] [3]),
        .O(\_T_2547[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hD0FFD0D0)) 
    \_T_2547[1]_i_1 
       (.I0(\req_tag_reg[0] ),
        .I1(\s2_req_tag_reg[6]_0 ),
        .I2(_T_2549[1]),
        .I3(\_T_2547[7]_i_3_n_0 ),
        .I4(\wb_reg_inst_reg[9]_0 ),
        .O(_T_2547[1]));
  (* SOFT_HLUTNM = "soft_lutpair1877" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \_T_2547[23]_i_3 
       (.I0(\_T_2547[31]_i_6_n_0 ),
        .I1(\reg_bp_0_control_tmatch_reg[1] [3]),
        .I2(\reg_bp_0_control_tmatch_reg[1] [4]),
        .O(\_T_2547[23]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1882" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \_T_2547[28]_i_3 
       (.I0(\reg_bp_0_control_tmatch_reg[1] [2]),
        .I1(\reg_bp_0_control_tmatch_reg[1] [1]),
        .I2(\reg_bp_0_control_tmatch_reg[1] [0]),
        .O(\_T_2547[28]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1883" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \_T_2547[29]_i_3 
       (.I0(\reg_bp_0_control_tmatch_reg[1] [2]),
        .I1(\reg_bp_0_control_tmatch_reg[1] [0]),
        .I2(\reg_bp_0_control_tmatch_reg[1] [1]),
        .O(\_T_2547[29]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hD0FFD0D0)) 
    \_T_2547[2]_i_1 
       (.I0(\req_tag_reg[1] ),
        .I1(\s2_req_tag_reg[6]_0 ),
        .I2(_T_2549[2]),
        .I3(\_T_2547[7]_i_3_n_0 ),
        .I4(\wb_reg_inst_reg[9]_1 ),
        .O(_T_2547[2]));
  (* SOFT_HLUTNM = "soft_lutpair1883" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \_T_2547[30]_i_3 
       (.I0(\reg_bp_0_control_tmatch_reg[1] [2]),
        .I1(\reg_bp_0_control_tmatch_reg[1] [1]),
        .I2(\reg_bp_0_control_tmatch_reg[1] [0]),
        .O(\_T_2547[30]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1876" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \_T_2547[31]_i_4 
       (.I0(\reg_bp_0_control_tmatch_reg[1] [4]),
        .I1(\_T_2547[31]_i_6_n_0 ),
        .I2(\reg_bp_0_control_tmatch_reg[1] [3]),
        .O(\_T_2547[31]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1882" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \_T_2547[31]_i_5 
       (.I0(\reg_bp_0_control_tmatch_reg[1] [2]),
        .I1(\reg_bp_0_control_tmatch_reg[1] [1]),
        .I2(\reg_bp_0_control_tmatch_reg[1] [0]),
        .O(\_T_2547[31]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h44440040)) 
    \_T_2547[31]_i_6 
       (.I0(wb_reg_replay_reg_0),
        .I1(wb_ctrl_wxd),
        .I2(wb_ctrl_mem),
        .I3(dcacheArb_io_requestor_1_resp_valid),
        .I4(wb_ctrl_div),
        .O(\_T_2547[31]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hD0FFD0D0)) 
    \_T_2547[3]_i_1 
       (.I0(\req_tag_reg[1]_0 ),
        .I1(\s2_req_tag_reg[6]_0 ),
        .I2(_T_2549[3]),
        .I3(\_T_2547[7]_i_3_n_0 ),
        .I4(\wb_reg_inst_reg[9]_2 ),
        .O(_T_2547[3]));
  LUT5 #(
    .INIT(32'hD0FFD0D0)) 
    \_T_2547[4]_i_1 
       (.I0(\req_tag_reg[1]_1 ),
        .I1(\s2_req_tag_reg[6]_0 ),
        .I2(_T_2549[4]),
        .I3(\_T_2547[7]_i_3_n_0 ),
        .I4(\_T_2547[28]_i_3_n_0 ),
        .O(_T_2547[4]));
  LUT5 #(
    .INIT(32'hD0FFD0D0)) 
    \_T_2547[5]_i_1 
       (.I0(\req_tag_reg[0]_0 ),
        .I1(\s2_req_tag_reg[6]_0 ),
        .I2(_T_2549[5]),
        .I3(\_T_2547[7]_i_3_n_0 ),
        .I4(\_T_2547[29]_i_3_n_0 ),
        .O(_T_2547[5]));
  LUT5 #(
    .INIT(32'hD0FFD0D0)) 
    \_T_2547[6]_i_1 
       (.I0(\req_tag_reg[1]_2 ),
        .I1(\s2_req_tag_reg[6]_0 ),
        .I2(_T_2549[6]),
        .I3(\_T_2547[7]_i_3_n_0 ),
        .I4(\_T_2547[30]_i_3_n_0 ),
        .O(_T_2547[6]));
  LUT5 #(
    .INIT(32'hD0FFD0D0)) 
    \_T_2547[7]_i_1 
       (.I0(\req_tag_reg[1]_3 ),
        .I1(\s2_req_tag_reg[6]_0 ),
        .I2(_T_2549[7]),
        .I3(\_T_2547[7]_i_3_n_0 ),
        .I4(\_T_2547[31]_i_5_n_0 ),
        .O(_T_2547[7]));
  (* SOFT_HLUTNM = "soft_lutpair1876" *) 
  LUT3 #(
    .INIT(8'hFD)) 
    \_T_2547[7]_i_3 
       (.I0(\_T_2547[31]_i_6_n_0 ),
        .I1(\reg_bp_0_control_tmatch_reg[1] [4]),
        .I2(\reg_bp_0_control_tmatch_reg[1] [3]),
        .O(\_T_2547[7]_i_3_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[10] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[10]),
        .Q(_T_2549[10]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[11] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[11]),
        .Q(_T_2549[11]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[12] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[12]),
        .Q(_T_2549[12]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[13] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[13]),
        .Q(_T_2549[13]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[14] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[14]),
        .Q(_T_2549[14]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[15] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[15]),
        .Q(_T_2549[15]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[16] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[16]),
        .Q(\_T_2547_reg[16]_0 ),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[17] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[17]),
        .Q(_T_2549[17]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[18] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[18]),
        .Q(_T_2549[18]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[19] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[19]),
        .Q(_T_2549[19]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[1] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[1]),
        .Q(_T_2549[1]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[20] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[20]),
        .Q(_T_2549[20]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[21] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[21]),
        .Q(_T_2549[21]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[22] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[22]),
        .Q(_T_2549[22]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[23] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[23]),
        .Q(_T_2549[23]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[24] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[24]),
        .Q(_T_2549[24]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[25] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[25]),
        .Q(_T_2549[25]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[26] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[26]),
        .Q(_T_2549[26]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[27] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[27]),
        .Q(_T_2549[27]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[28] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[28]),
        .Q(_T_2549[28]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[29] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[29]),
        .Q(_T_2549[29]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[2] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[2]),
        .Q(_T_2549[2]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[30] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[30]),
        .Q(_T_2549[30]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[31] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[31]),
        .Q(_T_2549[31]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[3] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[3]),
        .Q(_T_2549[3]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[4] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[4]),
        .Q(_T_2549[4]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[5] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[5]),
        .Q(_T_2549[5]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[6] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[6]),
        .Q(_T_2549[6]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[7] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[7]),
        .Q(_T_2549[7]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[8] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[8]),
        .Q(_T_2549[8]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \_T_2547_reg[9] 
       (.C(host_clk),
        .CE(E),
        .D(_T_2547[9]),
        .Q(_T_2549[9]),
        .R(target_reset));
  (* SOFT_HLUTNM = "soft_lutpair1879" *) 
  LUT3 #(
    .INIT(8'hBA)) 
    \_T_389[7]_i_1 
       (.I0(target_reset),
        .I1(\valid_reg[3]_1 ),
        .I2(frontend_io_cpu_sfence_valid),
        .O(\_T_389_reg[7] ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[0]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[0]),
        .I1(\bypass_mux_1[0]_i_2_n_0 ),
        .I2(\bypass_mux_1[0]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[0]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[0]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(\bypass_mux_1_reg[0]_0 ),
        .I2(alu_io_in2[0]),
        .I3(\bypass_mux_1[0]_i_4_n_0 ),
        .I4(core__160_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0FFF0FFFFFBBFFFF)) 
    \bypass_mux_1[0]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(\bypass_mux_1[0]_i_5_n_0 ),
        .I2(\bypass_mux_1[0]_i_6_n_0 ),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .I5(Q),
        .O(\bypass_mux_1[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[0]_i_4 
       (.I0(alu_io_in2[0]),
        .I1(\bypass_mux_1_reg[0]_0 ),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[0]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1832" *) 
  LUT4 #(
    .INIT(16'hCDC8)) 
    \bypass_mux_1[0]_i_5 
       (.I0(alu_io_in2[0]),
        .I1(_T_121),
        .I2(alu_io_in2[1]),
        .I3(\bypass_mux_1_reg[1]_1 ),
        .O(\bypass_mux_1[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hC5AC)) 
    \bypass_mux_1[0]_i_6 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(\ex_reg_pc_reg[39]_1 ),
        .I2(alu_io_in2[62]),
        .I3(alu_io_in1[62]),
        .O(\bypass_mux_1[0]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[10]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[10]),
        .I1(\bypass_mux_1[10]_i_2_n_0 ),
        .I2(\bypass_mux_1[10]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[10]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[10]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[9]),
        .I2(alu_io_in2[9]),
        .I3(\bypass_mux_1[10]_i_4_n_0 ),
        .I4(core__150_i_4_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[10]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_10),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[10]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[10]_i_4 
       (.I0(alu_io_in2[9]),
        .I1(alu_io_in1[9]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[10]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[11]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[11]),
        .I1(\bypass_mux_1[11]_i_3_n_0 ),
        .I2(\bypass_mux_1[11]_i_4_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[11]));
  LUT5 #(
    .INIT(32'h002A2A2A)) 
    \bypass_mux_1[11]_i_3 
       (.I0(\bypass_mux_1[11]_i_5_n_0 ),
        .I1(\ex_ctrl_alu_fn_reg[3]_0 ),
        .I2(\alu/_T_198 ),
        .I3(core__149_i_5_n_0),
        .I4(\alu/_T_55 ),
        .O(\bypass_mux_1[11]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[11]_i_4 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_9),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[11]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    \bypass_mux_1[11]_i_5 
       (.I0(alu_io_in2[10]),
        .I1(alu_io_in1[10]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1[11]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[12]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[12]),
        .I1(\bypass_mux_1[12]_i_2_n_0 ),
        .I2(\bypass_mux_1[12]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[12]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[12]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[11]),
        .I2(alu_io_in2[11]),
        .I3(\bypass_mux_1[12]_i_4_n_0 ),
        .I4(core__148_i_4_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[12]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[12]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_8),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[12]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[12]_i_4 
       (.I0(alu_io_in2[11]),
        .I1(alu_io_in1[11]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[12]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[13]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[13]),
        .I1(\bypass_mux_1[13]_i_2_n_0 ),
        .I2(\bypass_mux_1[13]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[13]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[13]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[12]),
        .I2(alu_io_in2[12]),
        .I3(\bypass_mux_1[13]_i_4_n_0 ),
        .I4(core__147_i_4_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[13]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[13]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_7),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[13]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[13]_i_4 
       (.I0(alu_io_in2[12]),
        .I1(alu_io_in1[12]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[13]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[14]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[14]),
        .I1(\bypass_mux_1[14]_i_2_n_0 ),
        .I2(\bypass_mux_1[14]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[14]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[14]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[13]),
        .I2(alu_io_in2[13]),
        .I3(\bypass_mux_1[14]_i_4_n_0 ),
        .I4(core__146_i_4_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[14]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_6),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[14]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[14]_i_4 
       (.I0(alu_io_in2[13]),
        .I1(alu_io_in1[13]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[14]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[15]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[15]),
        .I1(\bypass_mux_1[15]_i_3_n_0 ),
        .I2(\bypass_mux_1[15]_i_4_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[15]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[15]_i_3 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[14]),
        .I2(alu_io_in2[14]),
        .I3(\bypass_mux_1[15]_i_5_n_0 ),
        .I4(core__145_i_5_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[15]_i_4 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_5),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[15]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[15]_i_5 
       (.I0(alu_io_in2[14]),
        .I1(alu_io_in1[14]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[15]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[16]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[16]),
        .I1(\bypass_mux_1[16]_i_2_n_0 ),
        .I2(\bypass_mux_1[16]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[16]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[16]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[15]),
        .I2(alu_io_in2[15]),
        .I3(\bypass_mux_1[16]_i_4_n_0 ),
        .I4(core__144_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[16]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[16]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_4),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[16]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[16]_i_4 
       (.I0(alu_io_in2[15]),
        .I1(alu_io_in1[15]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[16]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[17]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[17]),
        .I1(\bypass_mux_1[17]_i_2_n_0 ),
        .I2(\bypass_mux_1[17]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[17]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[17]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[16]),
        .I2(alu_io_in2[16]),
        .I3(\bypass_mux_1[17]_i_4_n_0 ),
        .I4(core__143_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[17]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[17]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__143_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[17]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[17]_i_4 
       (.I0(alu_io_in2[16]),
        .I1(alu_io_in1[16]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[17]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[18]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[18]),
        .I1(\bypass_mux_1[18]_i_2_n_0 ),
        .I2(\bypass_mux_1[18]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[18]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[18]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[17]),
        .I2(alu_io_in2[17]),
        .I3(\bypass_mux_1[18]_i_4_n_0 ),
        .I4(core__142_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[18]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__142_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[18]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[18]_i_4 
       (.I0(alu_io_in2[17]),
        .I1(alu_io_in1[17]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[18]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[19]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[19]),
        .I1(\bypass_mux_1[19]_i_3_n_0 ),
        .I2(\bypass_mux_1[19]_i_4_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[19]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[19]_i_3 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[18]),
        .I2(alu_io_in2[18]),
        .I3(\bypass_mux_1[19]_i_5_n_0 ),
        .I4(core__141_i_4_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[19]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[19]_i_4 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__141_i_6_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[19]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[19]_i_5 
       (.I0(alu_io_in2[18]),
        .I1(alu_io_in1[18]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[19]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAAAACFFF)) 
    \bypass_mux_1[1]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[1]),
        .I1(\bypass_mux_1[1]_i_2_n_0 ),
        .I2(\bypass_mux_1[1]_i_3_n_0 ),
        .I3(\bypass_mux_1[1]_i_4_n_0 ),
        .I4(_T_217),
        .O(alu_io_out[1]));
  LUT6 #(
    .INIT(64'hFFFF8A808A808A80)) 
    \bypass_mux_1[1]_i_2 
       (.I0(\alu/_T_55 ),
        .I1(core__159_i_4_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__159_i_3_n_0),
        .I4(\alu/_T_198 ),
        .I5(\ex_ctrl_alu_fn_reg[3]_1 ),
        .O(\bypass_mux_1[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    \bypass_mux_1[1]_i_3 
       (.I0(alu_io_in2[1]),
        .I1(alu_io_in1[0]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[1]_i_4 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(\bypass_mux_1[1]_i_5_n_0 ),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[1]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1832" *) 
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    \bypass_mux_1[1]_i_5 
       (.I0(\bypass_mux_1_reg[1]_1 ),
        .I1(alu_io_in2[0]),
        .I2(_T_121),
        .I3(alu_io_in2[1]),
        .I4(\bypass_mux_1_reg[1]_2 ),
        .O(\bypass_mux_1[1]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[20]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[20]),
        .I1(\bypass_mux_1[20]_i_2_n_0 ),
        .I2(\bypass_mux_1[20]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[20]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[20]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[19]),
        .I2(alu_io_in2[19]),
        .I3(\bypass_mux_1[20]_i_4_n_0 ),
        .I4(core__140_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[20]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[20]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__140_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[20]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[20]_i_4 
       (.I0(alu_io_in2[19]),
        .I1(alu_io_in1[19]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[20]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[21]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[21]),
        .I1(\bypass_mux_1[21]_i_2_n_0 ),
        .I2(\bypass_mux_1[21]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[21]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[21]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[20]),
        .I2(alu_io_in2[20]),
        .I3(\bypass_mux_1[21]_i_4_n_0 ),
        .I4(core__139_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[21]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[21]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__139_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[21]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[21]_i_4 
       (.I0(alu_io_in2[20]),
        .I1(alu_io_in1[20]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[21]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[22]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[22]),
        .I1(\bypass_mux_1[22]_i_2_n_0 ),
        .I2(\bypass_mux_1[22]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[22]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[22]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[21]),
        .I2(alu_io_in2[21]),
        .I3(\bypass_mux_1[22]_i_4_n_0 ),
        .I4(core__138_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[22]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[22]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__138_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[22]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[22]_i_4 
       (.I0(alu_io_in2[21]),
        .I1(alu_io_in1[21]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[22]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[23]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[23]),
        .I1(\bypass_mux_1[23]_i_3_n_0 ),
        .I2(\bypass_mux_1[23]_i_4_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[23]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[23]_i_3 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[22]),
        .I2(alu_io_in2[22]),
        .I3(\bypass_mux_1[23]_i_5_n_0 ),
        .I4(core__137_i_4_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[23]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[23]_i_4 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__137_i_6_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[23]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[23]_i_5 
       (.I0(alu_io_in2[22]),
        .I1(alu_io_in1[22]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[23]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[24]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[24]),
        .I1(\bypass_mux_1[24]_i_2_n_0 ),
        .I2(\bypass_mux_1[24]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[24]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[24]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[23]),
        .I2(alu_io_in2[23]),
        .I3(\bypass_mux_1[24]_i_4_n_0 ),
        .I4(core__136_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[24]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[24]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__136_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[24]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[24]_i_4 
       (.I0(alu_io_in2[23]),
        .I1(alu_io_in1[23]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[24]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[25]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[25]),
        .I1(\bypass_mux_1[25]_i_2_n_0 ),
        .I2(\bypass_mux_1[25]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[25]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[25]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[24]),
        .I2(alu_io_in2[24]),
        .I3(\bypass_mux_1[25]_i_4_n_0 ),
        .I4(core__135_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[25]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[25]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__135_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[25]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[25]_i_4 
       (.I0(alu_io_in2[24]),
        .I1(alu_io_in1[24]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[25]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[26]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[26]),
        .I1(\bypass_mux_1[26]_i_2_n_0 ),
        .I2(\bypass_mux_1[26]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[26]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[26]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[25]),
        .I2(alu_io_in2[25]),
        .I3(\bypass_mux_1[26]_i_4_n_0 ),
        .I4(core__134_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[26]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[26]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__134_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[26]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[26]_i_4 
       (.I0(alu_io_in2[25]),
        .I1(alu_io_in1[25]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[26]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[27]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[27]),
        .I1(\bypass_mux_1[27]_i_3_n_0 ),
        .I2(\bypass_mux_1[27]_i_4_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[27]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[27]_i_3 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[26]),
        .I2(alu_io_in2[26]),
        .I3(\bypass_mux_1[27]_i_5_n_0 ),
        .I4(core__133_i_4_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[27]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[27]_i_4 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__133_i_6_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[27]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[27]_i_5 
       (.I0(alu_io_in2[26]),
        .I1(alu_io_in1[26]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[27]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[28]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[28]),
        .I1(\bypass_mux_1[28]_i_2_n_0 ),
        .I2(\bypass_mux_1[28]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[28]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[28]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[27]),
        .I2(alu_io_in2[27]),
        .I3(\bypass_mux_1[28]_i_4_n_0 ),
        .I4(core__132_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[28]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[28]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__132_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[28]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[28]_i_4 
       (.I0(alu_io_in2[27]),
        .I1(alu_io_in1[27]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[28]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[29]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[29]),
        .I1(\bypass_mux_1[29]_i_2_n_0 ),
        .I2(\bypass_mux_1[29]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[29]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[29]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[28]),
        .I2(alu_io_in2[28]),
        .I3(\bypass_mux_1[29]_i_4_n_0 ),
        .I4(core__131_i_3_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[29]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[29]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__131_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[29]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[29]_i_4 
       (.I0(alu_io_in2[28]),
        .I1(alu_io_in1[28]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[29]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAAACFFF)) 
    \bypass_mux_1[2]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[2]),
        .I1(\bypass_mux_1[2]_i_2_n_0 ),
        .I2(\bypass_mux_1[2]_i_3_n_0 ),
        .I3(\bypass_mux_1[2]_i_4_n_0 ),
        .I4(_T_217),
        .O(alu_io_out[2]));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    \bypass_mux_1[2]_i_2 
       (.I0(\alu/_T_55 ),
        .I1(core__158_i_3_n_0),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[1]),
        .I4(alu_io_in2[2]),
        .I5(Q),
        .O(\bypass_mux_1[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    \bypass_mux_1[2]_i_3 
       (.I0(alu_io_in2[2]),
        .I1(alu_io_in1[1]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[2]_i_4 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(\ex_ctrl_alu_fn_reg[3]_7 ),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[2]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[30]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[30]),
        .I1(\bypass_mux_1[30]_i_2_n_0 ),
        .I2(\bypass_mux_1[30]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[30]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[30]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[29]),
        .I2(alu_io_in2[29]),
        .I3(\bypass_mux_1[30]_i_4_n_0 ),
        .I4(ex_reg_rvc_reg_2),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[30]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[30]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_3),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[30]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[30]_i_4 
       (.I0(alu_io_in2[29]),
        .I1(alu_io_in1[29]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[30]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bypass_mux_1[31]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[31]),
        .I1(\bypass_mux_1_reg[32]_0 ),
        .I2(_T_217),
        .O(alu_io_out[31]));
  LUT6 #(
    .INIT(64'hAAAACCCCF0F0FF00)) 
    \bypass_mux_1[32]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[32]),
        .I1(dcacheArb_io_requestor_1_req_bits_addr[31]),
        .I2(\bypass_mux_1[32]_i_2_n_0 ),
        .I3(\bypass_mux_1_reg[32]_0 ),
        .I4(req_dw_reg),
        .I5(_T_217),
        .O(alu_io_out[32]));
  LUT5 #(
    .INIT(32'hEAAAFFFF)) 
    \bypass_mux_1[32]_i_2 
       (.I0(\bypass_mux_1[32]_i_3_n_0 ),
        .I1(alu_io_in2[31]),
        .I2(alu_io_in1[31]),
        .I3(\alu/_T_205 ),
        .I4(\bypass_mux_1[32]_i_4_n_0 ),
        .O(\bypass_mux_1[32]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    \bypass_mux_1[32]_i_3 
       (.I0(\alu/_T_55 ),
        .I1(core__161_i_6_n_0),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[31]),
        .I4(alu_io_in2[31]),
        .I5(Q),
        .O(\bypass_mux_1[32]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[32]_i_4 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__161_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[32]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAAACFFF)) 
    \bypass_mux_1[3]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[3]),
        .I1(\bypass_mux_1[3]_i_3_n_0 ),
        .I2(\bypass_mux_1[3]_i_4_n_0 ),
        .I3(\bypass_mux_1[3]_i_5_n_0 ),
        .I4(_T_217),
        .O(alu_io_out[3]));
  LUT6 #(
    .INIT(64'hFFFF8A808A808A80)) 
    \bypass_mux_1[3]_i_3 
       (.I0(\alu/_T_55 ),
        .I1(core__156_i_4_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__157_i_4_n_0),
        .I4(\alu/_T_198 ),
        .I5(\ex_ctrl_alu_fn_reg[3]_2 ),
        .O(\bypass_mux_1[3]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    \bypass_mux_1[3]_i_4 
       (.I0(alu_io_in2[3]),
        .I1(alu_io_in1[2]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1[3]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[3]_i_5 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(\ex_ctrl_alu_fn_reg[3]_6 ),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[3]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bypass_mux_1[3]_i_6 
       (.I0(div_n_240),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .O(\s1_req_addr_reg[3] ));
  LUT5 #(
    .INIT(32'hAAAACFFF)) 
    \bypass_mux_1[4]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[4]),
        .I1(\bypass_mux_1[4]_i_2_n_0 ),
        .I2(\bypass_mux_1[4]_i_3_n_0 ),
        .I3(\bypass_mux_1[4]_i_4_n_0 ),
        .I4(_T_217),
        .O(alu_io_out[4]));
  LUT6 #(
    .INIT(64'hFFFF8A808A808A80)) 
    \bypass_mux_1[4]_i_2 
       (.I0(\alu/_T_55 ),
        .I1(core__155_i_4_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__156_i_4_n_0),
        .I4(\alu/_T_198 ),
        .I5(\ex_ctrl_alu_fn_reg[3]_3 ),
        .O(\bypass_mux_1[4]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    \bypass_mux_1[4]_i_3 
       (.I0(alu_io_in2[4]),
        .I1(alu_io_in1[3]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1[4]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[4]_i_4 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_16),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[4]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAAACFFF)) 
    \bypass_mux_1[5]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[5]),
        .I1(\bypass_mux_1[5]_i_2_n_0 ),
        .I2(\bypass_mux_1[5]_i_3_n_0 ),
        .I3(\bypass_mux_1[5]_i_4_n_0 ),
        .I4(_T_217),
        .O(alu_io_out[5]));
  LUT6 #(
    .INIT(64'hFFFF8A808A808A80)) 
    \bypass_mux_1[5]_i_2 
       (.I0(\alu/_T_55 ),
        .I1(core__154_i_4_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__155_i_4_n_0),
        .I4(\alu/_T_198 ),
        .I5(\ex_ctrl_alu_fn_reg[3]_4 ),
        .O(\bypass_mux_1[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    \bypass_mux_1[5]_i_3 
       (.I0(alu_io_in2[5]),
        .I1(alu_io_in1[4]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1[5]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[5]_i_4 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_15),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFCCCFFFF)) 
    \bypass_mux_1[6]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[6]),
        .I1(\bypass_mux_1[6]_i_2_n_0 ),
        .I2(\alu/_T_206 [6]),
        .I3(\alu/_T_205 ),
        .I4(\bypass_mux_1[6]_i_4_n_0 ),
        .I5(_T_217),
        .O(alu_io_out[6]));
  LUT6 #(
    .INIT(64'hFFFF8A808A808A80)) 
    \bypass_mux_1[6]_i_2 
       (.I0(\alu/_T_55 ),
        .I1(core__154_i_5_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__154_i_4_n_0),
        .I4(\alu/_T_198 ),
        .I5(\ex_reg_inst_reg[26]_0 ),
        .O(\bypass_mux_1[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h08080808AA080808)) 
    \bypass_mux_1[6]_i_3 
       (.I0(alu_io_in1[5]),
        .I1(\mem_reg_inst_reg[31]_0 [5]),
        .I2(\bypass_mux_1_reg[6]_0 ),
        .I3(\divisor_reg[57] [1]),
        .I4(ex_ctrl_sel_alu2[1]),
        .I5(ex_ctrl_sel_alu2[0]),
        .O(\alu/_T_206 [6]));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[6]_i_4 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_14),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFCCCFFFF)) 
    \bypass_mux_1[7]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[7]),
        .I1(\bypass_mux_1[7]_i_3_n_0 ),
        .I2(\alu/_T_206 [7]),
        .I3(\alu/_T_205 ),
        .I4(\bypass_mux_1[7]_i_6_n_0 ),
        .I5(_T_217),
        .O(alu_io_out[7]));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    \bypass_mux_1[7]_i_3 
       (.I0(\alu/_T_55 ),
        .I1(core__153_i_5_n_0),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[6]),
        .I4(alu_io_in2[6]),
        .I5(Q),
        .O(\bypass_mux_1[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h08080808AA080808)) 
    \bypass_mux_1[7]_i_4 
       (.I0(alu_io_in1[6]),
        .I1(\mem_reg_inst_reg[31]_0 [6]),
        .I2(\bypass_mux_1_reg[6]_0 ),
        .I3(\divisor_reg[57] [2]),
        .I4(ex_ctrl_sel_alu2[1]),
        .I5(ex_ctrl_sel_alu2[0]),
        .O(\alu/_T_206 [7]));
  LUT3 #(
    .INIT(8'h08)) 
    \bypass_mux_1[7]_i_5 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[2]),
        .I2(Q),
        .O(\alu/_T_205 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[7]_i_6 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_13),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[7]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[8]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[8]),
        .I1(\bypass_mux_1[8]_i_2_n_0 ),
        .I2(\bypass_mux_1[8]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[8]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[8]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[7]),
        .I2(alu_io_in2[7]),
        .I3(\bypass_mux_1[8]_i_4_n_0 ),
        .I4(core__152_i_4_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[8]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[8]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_12),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[8]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[8]_i_4 
       (.I0(alu_io_in2[7]),
        .I1(alu_io_in1[7]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[8]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hAA3F)) 
    \bypass_mux_1[9]_i_1 
       (.I0(dcacheArb_io_requestor_1_req_bits_addr[9]),
        .I1(\bypass_mux_1[9]_i_2_n_0 ),
        .I2(\bypass_mux_1[9]_i_3_n_0 ),
        .I3(_T_217),
        .O(alu_io_out[9]));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \bypass_mux_1[9]_i_2 
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[8]),
        .I2(alu_io_in2[8]),
        .I3(\bypass_mux_1[9]_i_4_n_0 ),
        .I4(core__151_i_4_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1[9]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \bypass_mux_1[9]_i_3 
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_11),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1[9]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    \bypass_mux_1[9]_i_4 
       (.I0(alu_io_in2[8]),
        .I1(alu_io_in1[8]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(\bypass_mux_1[9]_i_4_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[0] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[0]),
        .Q(\bypass_mux_1_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[10] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[10]),
        .Q(\bypass_mux_1_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[11] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[11]),
        .Q(\bypass_mux_1_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[12] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[12]),
        .Q(\bypass_mux_1_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[13] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[13]),
        .Q(\bypass_mux_1_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[14] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[14]),
        .Q(\bypass_mux_1_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[15] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[15]),
        .Q(\bypass_mux_1_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[16] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[16]),
        .Q(\bypass_mux_1_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[17] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[17]),
        .Q(\bypass_mux_1_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[18] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[18]),
        .Q(\bypass_mux_1_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[19] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[19]),
        .Q(\bypass_mux_1_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[1] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[1]),
        .Q(\mem_reg_rs2_reg[3]_1 [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[20] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[20]),
        .Q(\bypass_mux_1_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[21] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[21]),
        .Q(\bypass_mux_1_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[22] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[22]),
        .Q(\bypass_mux_1_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[23] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[23]),
        .Q(\bypass_mux_1_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[24] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[24]),
        .Q(\bypass_mux_1_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[25] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[25]),
        .Q(\bypass_mux_1_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[26] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[26]),
        .Q(\bypass_mux_1_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[27] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[27]),
        .Q(\bypass_mux_1_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[28] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[28]),
        .Q(\bypass_mux_1_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[29] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[29]),
        .Q(\bypass_mux_1_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[2] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[2]),
        .Q(\bypass_mux_1_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[30] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[30]),
        .Q(\bypass_mux_1_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[31] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[31]),
        .Q(\bypass_mux_1_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[32] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[32]),
        .Q(\bypass_mux_1_reg_n_0_[32] ),
        .R(\<const0> ));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[33] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_32),
        .Q(\bypass_mux_1_reg_n_0_[33] ),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[34] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_31),
        .Q(\bypass_mux_1_reg_n_0_[34] ),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[35] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_30),
        .Q(\bypass_mux_1_reg_n_0_[35] ),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[36] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_29),
        .Q(\bypass_mux_1_reg_n_0_[36] ),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[37] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_28),
        .Q(\bypass_mux_1_reg_n_0_[37] ),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[38] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_27),
        .Q(\bypass_mux_2_reg[38]_0 ),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[39] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_26),
        .Q(_T_2177[0]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[3] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[3]),
        .Q(\mem_reg_rs2_reg[3]_1 [1]),
        .R(\<const0> ));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[40] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_25),
        .Q(_T_2177[1]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[41] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_24),
        .Q(_T_2177[2]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[42] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_23),
        .Q(_T_2177[3]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[43] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_22),
        .Q(_T_2177[4]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[44] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_21),
        .Q(_T_2177[5]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[45] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_20),
        .Q(_T_2177[6]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[46] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_19),
        .Q(_T_2177[7]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[47] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_18),
        .Q(_T_2177[8]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[48] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_17),
        .Q(_T_2177[9]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[49] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_16),
        .Q(_T_2177[10]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[4] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[4]),
        .Q(\bypass_mux_1_reg_n_0_[4] ),
        .R(\<const0> ));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[50] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_15),
        .Q(_T_2177[11]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[51] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_14),
        .Q(_T_2177[12]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[52] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_13),
        .Q(_T_2177[13]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[53] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_12),
        .Q(_T_2177[14]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[54] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_11),
        .Q(_T_2177[15]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[55] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_10),
        .Q(_T_2177[16]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[56] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_9),
        .Q(_T_2177[17]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[57] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_8),
        .Q(_T_2177[18]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[58] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_7),
        .Q(_T_2177[19]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[59] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_6),
        .Q(_T_2177[20]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[5] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[5]),
        .Q(\bypass_mux_1_reg_n_0_[5] ),
        .R(\<const0> ));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[60] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_5),
        .Q(_T_2177[21]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[61] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_4),
        .Q(_T_2177[22]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[62] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_3),
        .Q(_T_2177[23]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDSE #(
    .INIT(1'b1)) 
    \bypass_mux_1_reg[63] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_alu_dw_reg_2),
        .Q(_T_2177[24]),
        .S(ex_ctrl_alu_dw_reg_1));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[6] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[6]),
        .Q(\bypass_mux_1_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[7] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[7]),
        .Q(\bypass_mux_1_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[8] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[8]),
        .Q(\bypass_mux_1_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_1_reg[9] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_out[9]),
        .Q(\bypass_mux_1_reg_n_0_[9] ),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'hA8)) 
    \bypass_mux_2[31]_i_3 
       (.I0(\wb_reg_inst_reg[31]_0 [24]),
        .I1(\bypass_mux_2_reg[35]_0 ),
        .I2(mem_ctrl_jal),
        .O(\bypass_mux_2_reg[31]_0 [3]));
  LUT3 #(
    .INIT(8'h1F)) 
    \bypass_mux_2[35]_i_3 
       (.I0(mem_ctrl_jal),
        .I1(\bypass_mux_2_reg[35]_0 ),
        .I2(\wb_reg_inst_reg[31]_0 [24]),
        .O(\wb_reg_pc_reg[34]_0 [0]));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[0] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[0]),
        .Q(\mem_reg_rs2_reg[0]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[10] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[10]),
        .Q(\reg_mtvec_reg[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[11] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[11]),
        .Q(\reg_mtvec_reg[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[12] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[12]),
        .Q(\reg_mtvec_reg[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[13] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[13]),
        .Q(\reg_mtvec_reg[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[14] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[14]),
        .Q(\reg_mtvec_reg[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[15] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[15]),
        .Q(\reg_mtvec_reg[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[16] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[16]),
        .Q(\reg_mtvec_reg[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[17] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[17]),
        .Q(\reg_mtvec_reg[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[18] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[18]),
        .Q(\reg_mtvec_reg[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[19] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[19]),
        .Q(\reg_mtvec_reg[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[1] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[1]),
        .Q(\mem_reg_rs2_reg[1]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[20] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[20]),
        .Q(\reg_mtvec_reg[20]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[21] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[21]),
        .Q(\reg_mtvec_reg[21]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[22] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[22]),
        .Q(\reg_mtvec_reg[22]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[23] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[23]),
        .Q(\reg_mtvec_reg[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[24] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[24]),
        .Q(\reg_mtvec_reg[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[25] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[25]),
        .Q(\reg_mtvec_reg[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[26] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[26]),
        .Q(\reg_mtvec_reg[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[27] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[27]),
        .Q(\reg_mtvec_reg[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[28] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[28]),
        .Q(\reg_mtvec_reg[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[29] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[29]),
        .Q(\reg_mtvec_reg[29]_7 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[2] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[2]),
        .Q(\mem_reg_rs2_reg[2]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[30] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[30]),
        .Q(\reg_mtvec_reg[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[31] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[31]),
        .Q(\reg_mtvec_reg[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[32] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[32]),
        .Q(\reg_stvec_reg[32] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[33] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[33]),
        .Q(\reg_stvec_reg[33] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[34] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[34]),
        .Q(\reg_stvec_reg[34] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[35] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[35]),
        .Q(\reg_stvec_reg[35] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[36] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[36]),
        .Q(\reg_stvec_reg[36] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[37] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[37]),
        .Q(\reg_stvec_reg[37] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[38] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[38]),
        .Q(\reg_stvec_reg[38] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[39] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[39]),
        .Q(\reg_sscratch_reg[62] [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[3] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[3]),
        .Q(\mem_reg_rs2_reg[3]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[40] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[40]),
        .Q(\reg_sscratch_reg[62] [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[41] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[41]),
        .Q(\reg_sscratch_reg[62] [2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[42] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[42]),
        .Q(\reg_sscratch_reg[62] [3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[43] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[43]),
        .Q(\reg_sscratch_reg[62] [4]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[44] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[44]),
        .Q(\reg_sscratch_reg[62] [5]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[45] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[45]),
        .Q(\reg_sscratch_reg[62] [6]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[46] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[46]),
        .Q(\reg_sscratch_reg[62] [7]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[47] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[47]),
        .Q(\reg_sscratch_reg[62] [8]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[48] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[48]),
        .Q(\reg_sscratch_reg[62] [9]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[49] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[49]),
        .Q(\reg_sscratch_reg[62] [10]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[4] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[4]),
        .Q(\mem_reg_rs2_reg[4]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[50] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[50]),
        .Q(\reg_sscratch_reg[62] [11]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[51] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[51]),
        .Q(\reg_sscratch_reg[62] [12]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[52] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[52]),
        .Q(\reg_sscratch_reg[62] [13]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[53] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[53]),
        .Q(\reg_sscratch_reg[62] [14]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[54] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[54]),
        .Q(\reg_sscratch_reg[62] [15]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[55] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[55]),
        .Q(\reg_sscratch_reg[62] [16]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[56] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[56]),
        .Q(\reg_sscratch_reg[62] [17]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[57] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[57]),
        .Q(\reg_sscratch_reg[62] [18]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[58] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[58]),
        .Q(\reg_sscratch_reg[62] [19]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[59] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[59]),
        .Q(\reg_sscratch_reg[62] [20]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[5] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[5]),
        .Q(\mem_reg_rs2_reg[5]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[60] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[60]),
        .Q(\reg_sscratch_reg[62] [21]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[61] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[61]),
        .Q(\reg_sscratch_reg[62] [22]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[62] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[62]),
        .Q(\reg_sscratch_reg[62] [23]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[63] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[63]),
        .Q(_T_2518),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[6] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[6]),
        .Q(\mem_reg_rs2_reg[6]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[7] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[7]),
        .Q(\mem_reg_rs2_reg[7]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[8] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[8]),
        .Q(\reg_mtvec_reg[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \bypass_mux_2_reg[9] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_int_wdata[9]),
        .Q(reg_mip_seip_reg_0),
        .R(\<const0> ));
  LUT5 #(
    .INIT(32'h00000040)) 
    core__115_i_1
       (.I0(core__115_i_2_n_0),
        .I1(wb_reg_valid),
        .I2(\reg_sscratch_reg[59] [2]),
        .I3(\reg_sscratch_reg[59] [1]),
        .I4(\reg_sscratch_reg[59] [0]),
        .O(reg_debug_reg));
  (* SOFT_HLUTNM = "soft_lutpair1864" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    core__115_i_2
       (.I0(\reg_bp_0_control_tmatch_reg[1] [7]),
        .I1(\reg_bp_0_control_tmatch_reg[1] [6]),
        .I2(\reg_bp_0_control_tmatch_reg[1] [5]),
        .O(core__115_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1783" *) 
  LUT5 #(
    .INIT(32'h00000008)) 
    core__116_i_10
       (.I0(wb_reg_valid),
        .I1(\reg_sscratch_reg[59] [2]),
        .I2(\reg_sscratch_reg[59] [1]),
        .I3(\reg_sscratch_reg[59] [0]),
        .I4(core__116_i_11_n_0),
        .O(core__116_i_10_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1864" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    core__116_i_11
       (.I0(\reg_bp_0_control_tmatch_reg[1] [7]),
        .I1(\reg_bp_0_control_tmatch_reg[1] [5]),
        .I2(\reg_bp_0_control_tmatch_reg[1] [6]),
        .O(core__116_i_11_n_0));
  LUT4 #(
    .INIT(16'h0041)) 
    core__130_i_1
       (.I0(ex_ctrl_alu_fn[0]),
        .I1(ex_ctrl_alu_fn[1]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .O(_T_217));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__130_i_2
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(ex_reg_rvc_reg_2),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[33]_1 ));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__130_i_3
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[32]),
        .I2(alu_io_in2[32]),
        .I3(core__130_i_5_n_0),
        .I4(ex_reg_rvc_reg_3),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[33]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__130_i_5
       (.I0(alu_io_in2[32]),
        .I1(alu_io_in1[32]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__130_i_5_n_0));
  LUT4 #(
    .INIT(16'h1800)) 
    core__130_i_6
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(Q),
        .I2(ex_ctrl_alu_fn[2]),
        .I3(ex_ctrl_alu_fn[0]),
        .O(\alu/_T_55 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__131_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__131_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[34]_1 ));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__131_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[33]),
        .I2(alu_io_in2[33]),
        .I3(core__131_i_4_n_0),
        .I4(core__131_i_5_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[34]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__131_i_3
       (.I0(\bypass_mux_1_reg[34]_2 ),
        .I1(\ex_reg_inst_reg[10]_4 ),
        .I2(alu_io_in2[0]),
        .I3(\bypass_mux_1_reg[35]_2 ),
        .I4(alu_io_in2[1]),
        .I5(\ex_reg_inst_reg[10]_3 ),
        .O(core__131_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__131_i_4
       (.I0(alu_io_in2[33]),
        .I1(alu_io_in1[33]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__131_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__131_i_5
       (.I0(\ex_reg_inst_reg[10]_5 ),
        .I1(\bypass_mux_1_reg[29]_1 ),
        .I2(alu_io_in2[0]),
        .I3(\ex_reg_inst_reg[10]_6 ),
        .I4(alu_io_in2[1]),
        .I5(\bypass_mux_1_reg[29]_0 ),
        .O(core__131_i_5_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__132_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__132_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[35]_1 ));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__132_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[34]),
        .I2(alu_io_in2[34]),
        .I3(core__132_i_4_n_0),
        .I4(core__132_i_5_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[35]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__132_i_3
       (.I0(\bypass_mux_1_reg[35]_2 ),
        .I1(\ex_reg_inst_reg[10]_3 ),
        .I2(alu_io_in2[0]),
        .I3(\ex_reg_inst_reg[10]_4 ),
        .I4(alu_io_in2[1]),
        .I5(\ex_reg_inst_reg[10]_2 ),
        .O(core__132_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__132_i_4
       (.I0(alu_io_in2[34]),
        .I1(alu_io_in1[34]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__132_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__132_i_5
       (.I0(\ex_reg_inst_reg[10]_7 ),
        .I1(\ex_reg_inst_reg[10]_6 ),
        .I2(alu_io_in2[0]),
        .I3(\ex_reg_inst_reg[10]_5 ),
        .I4(alu_io_in2[1]),
        .I5(\bypass_mux_1_reg[29]_1 ),
        .O(core__132_i_5_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__133_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__133_i_4_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[36]_1 ));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__133_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[35]),
        .I2(alu_io_in2[35]),
        .I3(core__133_i_5_n_0),
        .I4(core__133_i_6_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[36]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__133_i_4
       (.I0(\ex_reg_inst_reg[10]_4 ),
        .I1(\ex_reg_inst_reg[10]_2 ),
        .I2(alu_io_in2[0]),
        .I3(\ex_reg_inst_reg[10]_3 ),
        .I4(alu_io_in2[1]),
        .I5(\ex_reg_inst_reg[10]_1 ),
        .O(core__133_i_4_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__133_i_5
       (.I0(alu_io_in2[35]),
        .I1(alu_io_in1[35]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__133_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__133_i_6
       (.I0(\ex_ctrl_alu_fn_reg[3]_5 ),
        .I1(\ex_reg_inst_reg[10]_5 ),
        .I2(alu_io_in2[0]),
        .I3(\ex_reg_inst_reg[10]_7 ),
        .I4(alu_io_in2[1]),
        .I5(\ex_reg_inst_reg[10]_6 ),
        .O(core__133_i_6_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__134_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__134_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[37]_1 ));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__134_i_10
       (.I0(\alu/shin [58]),
        .I1(shamt),
        .I2(alu_io_in1[25]),
        .I3(core__134_i_11_n_0),
        .I4(\alu/_T_55 ),
        .O(core__134_i_10_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1816" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__134_i_11
       (.I0(alu_io_in1[36]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__134_i_11_n_0));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__134_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[36]),
        .I2(alu_io_in2[36]),
        .I3(core__134_i_4_n_0),
        .I4(core__134_i_5_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[37]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__134_i_3
       (.I0(\ex_reg_inst_reg[10]_3 ),
        .I1(\ex_reg_inst_reg[10]_1 ),
        .I2(alu_io_in2[0]),
        .I3(\ex_reg_inst_reg[10]_2 ),
        .I4(alu_io_in2[1]),
        .I5(core__134_i_6_n_0),
        .O(core__134_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__134_i_4
       (.I0(alu_io_in2[36]),
        .I1(alu_io_in1[36]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__134_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__134_i_5
       (.I0(core__134_i_7_n_0),
        .I1(\ex_reg_inst_reg[10]_7 ),
        .I2(alu_io_in2[0]),
        .I3(\ex_ctrl_alu_fn_reg[3]_5 ),
        .I4(alu_io_in2[1]),
        .I5(\ex_reg_inst_reg[10]_5 ),
        .O(core__134_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__134_i_6
       (.I0(\bypass_mux_1_reg[37]_2 ),
        .I1(\bypass_mux_1_reg[45]_2 ),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[41]_2 ),
        .I4(alu_io_in2[3]),
        .I5(core__134_i_8_n_0),
        .O(core__134_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1866" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__134_i_7
       (.I0(core__134_i_9_n_0),
        .I1(alu_io_in2[2]),
        .I2(\bypass_mux_1_reg[23]_0 ),
        .O(core__134_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__134_i_8
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [42]),
        .I3(alu_io_in2[4]),
        .I4(core__134_i_10_n_0),
        .O(core__134_i_8_n_0));
  LUT6 #(
    .INIT(64'hCDC8FFFFCDC80000)) 
    core__134_i_9
       (.I0(alu_io_in2[4]),
        .I1(_T_121),
        .I2(shamt),
        .I3(\alu/shin [52]),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[34]_3 ),
        .O(core__134_i_9_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__135_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__135_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[38]_1 ));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__135_i_10
       (.I0(\alu/shin [57]),
        .I1(shamt),
        .I2(alu_io_in1[24]),
        .I3(core__135_i_11_n_0),
        .I4(\alu/_T_55 ),
        .O(core__135_i_10_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1815" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__135_i_11
       (.I0(alu_io_in1[37]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__135_i_11_n_0));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__135_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[37]),
        .I2(alu_io_in2[37]),
        .I3(core__135_i_4_n_0),
        .I4(core__135_i_5_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[38]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__135_i_3
       (.I0(\ex_reg_inst_reg[10]_2 ),
        .I1(core__134_i_6_n_0),
        .I2(alu_io_in2[0]),
        .I3(\ex_reg_inst_reg[10]_1 ),
        .I4(alu_io_in2[1]),
        .I5(core__135_i_6_n_0),
        .O(core__135_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__135_i_4
       (.I0(alu_io_in2[37]),
        .I1(alu_io_in1[37]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__135_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__135_i_5
       (.I0(core__135_i_7_n_0),
        .I1(\ex_ctrl_alu_fn_reg[3]_5 ),
        .I2(alu_io_in2[0]),
        .I3(core__134_i_7_n_0),
        .I4(alu_io_in2[1]),
        .I5(\ex_reg_inst_reg[10]_7 ),
        .O(core__135_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__135_i_6
       (.I0(\bypass_mux_1_reg[38]_2 ),
        .I1(\bypass_mux_1_reg[46]_2 ),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[42]_2 ),
        .I4(alu_io_in2[3]),
        .I5(core__135_i_8_n_0),
        .O(core__135_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1874" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__135_i_7
       (.I0(core__135_i_9_n_0),
        .I1(alu_io_in2[2]),
        .I2(\bypass_mux_1_reg[22]_0 ),
        .O(core__135_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__135_i_8
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [41]),
        .I3(alu_io_in2[4]),
        .I4(core__135_i_10_n_0),
        .O(core__135_i_8_n_0));
  LUT6 #(
    .INIT(64'hCDC8FFFFCDC80000)) 
    core__135_i_9
       (.I0(alu_io_in2[4]),
        .I1(_T_121),
        .I2(shamt),
        .I3(\alu/shin [53]),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[33]_3 ),
        .O(core__135_i_9_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__136_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__136_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[39]_1 ));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__136_i_10
       (.I0(\alu/shin [56]),
        .I1(shamt),
        .I2(alu_io_in1[23]),
        .I3(core__136_i_11_n_0),
        .I4(\alu/_T_55 ),
        .O(core__136_i_10_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1809" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__136_i_11
       (.I0(alu_io_in1[38]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__136_i_11_n_0));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__136_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[38]),
        .I2(alu_io_in2[38]),
        .I3(core__136_i_4_n_0),
        .I4(core__136_i_5_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[39]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__136_i_3
       (.I0(\ex_reg_inst_reg[10]_1 ),
        .I1(core__135_i_6_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__134_i_6_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__136_i_6_n_0),
        .O(core__136_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__136_i_4
       (.I0(alu_io_in2[38]),
        .I1(alu_io_in1[38]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__136_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__136_i_5
       (.I0(core__136_i_7_n_0),
        .I1(core__134_i_7_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__135_i_7_n_0),
        .I4(alu_io_in2[1]),
        .I5(\ex_ctrl_alu_fn_reg[3]_5 ),
        .O(core__136_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__136_i_6
       (.I0(\bypass_mux_1_reg[39]_2 ),
        .I1(\bypass_mux_1_reg[47]_2 ),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[43]_2 ),
        .I4(alu_io_in2[3]),
        .I5(core__136_i_8_n_0),
        .O(core__136_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1875" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__136_i_7
       (.I0(core__136_i_9_n_0),
        .I1(alu_io_in2[2]),
        .I2(\bypass_mux_1_reg[21]_0 ),
        .O(core__136_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__136_i_8
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [40]),
        .I3(alu_io_in2[4]),
        .I4(core__136_i_10_n_0),
        .O(core__136_i_8_n_0));
  LUT6 #(
    .INIT(64'hCDC8FFFFCDC80000)) 
    core__136_i_9
       (.I0(alu_io_in2[4]),
        .I1(_T_121),
        .I2(shamt),
        .I3(\alu/shin [54]),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[29]_2 ),
        .O(core__136_i_9_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__137_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__137_i_4_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[40]_1 ));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__137_i_10
       (.I0(\alu/shin [55]),
        .I1(shamt),
        .I2(alu_io_in1[22]),
        .I3(core__137_i_11_n_0),
        .I4(\alu/_T_55 ),
        .O(core__137_i_10_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1812" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__137_i_11
       (.I0(alu_io_in1[39]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__137_i_11_n_0));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__137_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[39]),
        .I2(alu_io_in2[39]),
        .I3(core__137_i_5_n_0),
        .I4(core__137_i_6_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[40]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__137_i_4
       (.I0(core__134_i_6_n_0),
        .I1(core__136_i_6_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__135_i_6_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__137_i_7_n_0),
        .O(core__137_i_4_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__137_i_5
       (.I0(alu_io_in2[39]),
        .I1(alu_io_in1[39]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__137_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__137_i_6
       (.I0(core__137_i_8_n_0),
        .I1(core__135_i_7_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__136_i_7_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__134_i_7_n_0),
        .O(core__137_i_6_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__137_i_7
       (.I0(\bypass_mux_1_reg[40]_2 ),
        .I1(\bypass_mux_1_reg[48]_2 ),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[44]_2 ),
        .I4(alu_io_in2[3]),
        .I5(core__137_i_9_n_0),
        .O(core__137_i_7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1873" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__137_i_8
       (.I0(core__649_i_12_n_0),
        .I1(alu_io_in2[2]),
        .I2(\bypass_mux_1_reg[20]_0 ),
        .O(core__137_i_8_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__137_i_9
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [39]),
        .I3(alu_io_in2[4]),
        .I4(core__137_i_10_n_0),
        .O(core__137_i_9_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__138_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__138_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[41]_1 ));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__138_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[40]),
        .I2(alu_io_in2[40]),
        .I3(core__138_i_4_n_0),
        .I4(core__138_i_5_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[41]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__138_i_3
       (.I0(core__135_i_6_n_0),
        .I1(core__137_i_7_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__136_i_6_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__138_i_6_n_0),
        .O(core__138_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__138_i_4
       (.I0(alu_io_in2[40]),
        .I1(alu_io_in1[40]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__138_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__138_i_5
       (.I0(core__138_i_7_n_0),
        .I1(core__136_i_7_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__137_i_8_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__135_i_7_n_0),
        .O(core__138_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__138_i_6
       (.I0(\bypass_mux_1_reg[41]_2 ),
        .I1(core__134_i_8_n_0),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[45]_2 ),
        .I4(alu_io_in2[3]),
        .I5(core__138_i_8_n_0),
        .O(core__138_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1878" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__138_i_7
       (.I0(core__649_i_8_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__134_i_9_n_0),
        .O(core__138_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__138_i_8
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [38]),
        .I3(alu_io_in2[4]),
        .I4(core__154_i_9_n_0),
        .O(core__138_i_8_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__139_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__139_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[42]_1 ));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__139_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[41]),
        .I2(alu_io_in2[41]),
        .I3(core__139_i_4_n_0),
        .I4(core__139_i_5_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[42]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__139_i_3
       (.I0(core__136_i_6_n_0),
        .I1(core__138_i_6_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__137_i_7_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__139_i_6_n_0),
        .O(core__139_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__139_i_4
       (.I0(alu_io_in2[41]),
        .I1(alu_io_in1[41]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__139_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__139_i_5
       (.I0(core__139_i_7_n_0),
        .I1(core__137_i_8_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__138_i_7_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__136_i_7_n_0),
        .O(core__139_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__139_i_6
       (.I0(\bypass_mux_1_reg[42]_2 ),
        .I1(core__135_i_8_n_0),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[46]_2 ),
        .I4(alu_io_in2[3]),
        .I5(core__139_i_8_n_0),
        .O(core__139_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1874" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__139_i_7
       (.I0(core__649_i_10_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__135_i_9_n_0),
        .O(core__139_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__139_i_8
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [37]),
        .I3(alu_io_in2[4]),
        .I4(core__159_i_8_n_0),
        .O(core__139_i_8_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__140_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__140_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[43]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair1805" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__140_i_10
       (.I0(alu_io_in1[42]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__140_i_10_n_0));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__140_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[42]),
        .I2(alu_io_in2[42]),
        .I3(core__140_i_4_n_0),
        .I4(core__140_i_5_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[43]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__140_i_3
       (.I0(core__137_i_7_n_0),
        .I1(core__139_i_6_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__138_i_6_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__140_i_6_n_0),
        .O(core__140_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__140_i_4
       (.I0(alu_io_in2[42]),
        .I1(alu_io_in1[42]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__140_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__140_i_5
       (.I0(core__140_i_7_n_0),
        .I1(core__138_i_7_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__139_i_7_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__137_i_8_n_0),
        .O(core__140_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__140_i_6
       (.I0(\bypass_mux_1_reg[43]_2 ),
        .I1(core__136_i_8_n_0),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[47]_2 ),
        .I4(alu_io_in2[3]),
        .I5(core__140_i_8_n_0),
        .O(core__140_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1870" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__140_i_7
       (.I0(core__649_i_6_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__136_i_9_n_0),
        .O(core__140_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__140_i_8
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [36]),
        .I3(alu_io_in2[4]),
        .I4(core__140_i_9_n_0),
        .O(core__140_i_8_n_0));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__140_i_9
       (.I0(\alu/shin [52]),
        .I1(shamt),
        .I2(alu_io_in1[19]),
        .I3(core__140_i_10_n_0),
        .I4(\alu/_T_55 ),
        .O(core__140_i_9_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__141_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__141_i_4_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[44]_1 ));
  (* SOFT_HLUTNM = "soft_lutpair1808" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__141_i_10
       (.I0(alu_io_in1[43]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__141_i_10_n_0));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__141_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[43]),
        .I2(alu_io_in2[43]),
        .I3(core__141_i_5_n_0),
        .I4(core__141_i_6_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[44]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__141_i_4
       (.I0(core__138_i_6_n_0),
        .I1(core__140_i_6_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__139_i_6_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__141_i_7_n_0),
        .O(core__141_i_4_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__141_i_5
       (.I0(alu_io_in2[43]),
        .I1(alu_io_in1[43]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__141_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__141_i_6
       (.I0(\bypass_mux_1_reg[19]_0 ),
        .I1(core__139_i_7_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__140_i_7_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__138_i_7_n_0),
        .O(core__141_i_6_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__141_i_7
       (.I0(\bypass_mux_1_reg[44]_2 ),
        .I1(core__137_i_9_n_0),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[48]_2 ),
        .I4(alu_io_in2[3]),
        .I5(core__141_i_8_n_0),
        .O(core__141_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__141_i_8
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [35]),
        .I3(alu_io_in2[4]),
        .I4(core__141_i_9_n_0),
        .O(core__141_i_8_n_0));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__141_i_9
       (.I0(\alu/shin [51]),
        .I1(shamt),
        .I2(alu_io_in1[18]),
        .I3(core__141_i_10_n_0),
        .I4(\alu/_T_55 ),
        .O(core__141_i_9_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__142_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__142_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[45]_1 ));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__142_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[44]),
        .I2(alu_io_in2[44]),
        .I3(core__142_i_4_n_0),
        .I4(core__142_i_5_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[45]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__142_i_3
       (.I0(core__139_i_6_n_0),
        .I1(core__141_i_7_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__140_i_6_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__142_i_6_n_0),
        .O(core__142_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__142_i_4
       (.I0(alu_io_in2[44]),
        .I1(alu_io_in1[44]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__142_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__142_i_5
       (.I0(\bypass_mux_1_reg[18]_0 ),
        .I1(core__140_i_7_n_0),
        .I2(alu_io_in2[0]),
        .I3(\bypass_mux_1_reg[19]_0 ),
        .I4(alu_io_in2[1]),
        .I5(core__139_i_7_n_0),
        .O(core__142_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__142_i_6
       (.I0(\bypass_mux_1_reg[45]_2 ),
        .I1(core__138_i_8_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__134_i_8_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__142_i_7_n_0),
        .O(core__142_i_6_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__142_i_7
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [34]),
        .I3(alu_io_in2[4]),
        .I4(core__142_i_8_n_0),
        .O(core__142_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__142_i_8
       (.I0(\alu/shin [50]),
        .I1(shamt),
        .I2(alu_io_in1[17]),
        .I3(core__142_i_9_n_0),
        .I4(\alu/_T_55 ),
        .O(core__142_i_8_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1807" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__142_i_9
       (.I0(alu_io_in1[44]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__142_i_9_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__143_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__143_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[46]_1 ));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__143_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[45]),
        .I2(alu_io_in2[45]),
        .I3(core__143_i_4_n_0),
        .I4(core__143_i_5_n_0),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[46]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__143_i_3
       (.I0(core__140_i_6_n_0),
        .I1(core__142_i_6_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__141_i_7_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__143_i_6_n_0),
        .O(core__143_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__143_i_4
       (.I0(alu_io_in2[45]),
        .I1(alu_io_in1[45]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__143_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__143_i_5
       (.I0(\bypass_mux_1_reg[17]_0 ),
        .I1(\bypass_mux_1_reg[19]_0 ),
        .I2(alu_io_in2[0]),
        .I3(\bypass_mux_1_reg[18]_0 ),
        .I4(alu_io_in2[1]),
        .I5(core__140_i_7_n_0),
        .O(core__143_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__143_i_6
       (.I0(\bypass_mux_1_reg[46]_2 ),
        .I1(core__139_i_8_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__135_i_8_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__143_i_7_n_0),
        .O(core__143_i_6_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__143_i_7
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [33]),
        .I3(alu_io_in2[4]),
        .I4(core__159_i_10_n_0),
        .O(core__143_i_7_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__144_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__144_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[47]_1 ));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    core__144_i_2
       (.I0(\alu/_T_205 ),
        .I1(alu_io_in1[46]),
        .I2(alu_io_in2[46]),
        .I3(core__144_i_4_n_0),
        .I4(ex_reg_rvc_reg_4),
        .I5(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[47]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__144_i_3
       (.I0(core__141_i_7_n_0),
        .I1(core__143_i_6_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__142_i_6_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__144_i_5_n_0),
        .O(core__144_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFF9FF)) 
    core__144_i_4
       (.I0(alu_io_in2[46]),
        .I1(alu_io_in1[46]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[0]),
        .O(core__144_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__144_i_5
       (.I0(\bypass_mux_1_reg[47]_2 ),
        .I1(core__140_i_8_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__136_i_8_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__144_i_6_n_0),
        .O(core__144_i_5_n_0));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__144_i_6
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [32]),
        .I3(alu_io_in2[4]),
        .I4(core__144_i_7_n_0),
        .O(core__144_i_6_n_0));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__144_i_7
       (.I0(\alu/shin [48]),
        .I1(shamt),
        .I2(alu_io_in1[15]),
        .I3(core__144_i_8_n_0),
        .I4(\alu/_T_55 ),
        .O(core__144_i_7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1804" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__144_i_8
       (.I0(alu_io_in1[46]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__144_i_8_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__145_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__145_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[48]_1 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__145_i_2
       (.I0(alu_io_in2[47]),
        .I1(alu_io_in1[47]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[48]_3 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__145_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_5),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[47]),
        .I4(alu_io_in2[47]),
        .I5(Q),
        .O(\bypass_mux_1_reg[48]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__145_i_5
       (.I0(core__142_i_6_n_0),
        .I1(core__144_i_5_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__143_i_6_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__145_i_7_n_0),
        .O(core__145_i_5_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1802" *) 
  LUT3 #(
    .INIT(8'h04)) 
    core__145_i_6
       (.I0(ex_ctrl_alu_fn[0]),
        .I1(ex_ctrl_alu_fn[2]),
        .I2(Q),
        .O(\alu/_T_198 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__145_i_7
       (.I0(\bypass_mux_1_reg[48]_2 ),
        .I1(core__141_i_8_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__137_i_9_n_0),
        .I4(alu_io_in2[3]),
        .I5(ex_ctrl_alu_dw_reg_33),
        .O(core__145_i_7_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__146_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__146_i_4_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[49]_1 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__146_i_2
       (.I0(alu_io_in2[48]),
        .I1(alu_io_in1[48]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[49]_2 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__146_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_6),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[48]),
        .I4(alu_io_in2[48]),
        .I5(Q),
        .O(\bypass_mux_1_reg[49]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__146_i_4
       (.I0(core__143_i_6_n_0),
        .I1(core__145_i_7_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__144_i_5_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__146_i_5_n_0),
        .O(core__146_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__146_i_5
       (.I0(core__134_i_8_n_0),
        .I1(core__142_i_7_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__138_i_8_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__146_i_6_n_0),
        .O(core__146_i_5_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__146_i_6
       (.I0(core__644_i_12_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [46]),
        .I3(shamt),
        .I4(\alu/shin [14]),
        .O(core__146_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1785" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__146_i_7
       (.I0(alu_io_in1[13]),
        .I1(alu_io_in1[48]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [14]));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__147_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__147_i_4_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[50]_1 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__147_i_2
       (.I0(alu_io_in2[49]),
        .I1(alu_io_in1[49]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[50]_3 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__147_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_7),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[49]),
        .I4(alu_io_in2[49]),
        .I5(Q),
        .O(\bypass_mux_1_reg[50]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__147_i_4
       (.I0(core__144_i_5_n_0),
        .I1(core__146_i_5_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__145_i_7_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__147_i_5_n_0),
        .O(core__147_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__147_i_5
       (.I0(core__135_i_8_n_0),
        .I1(core__143_i_7_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__139_i_8_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__147_i_6_n_0),
        .O(core__147_i_5_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__147_i_6
       (.I0(core__643_i_12_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [45]),
        .I3(shamt),
        .I4(\alu/shin [13]),
        .O(core__147_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1801" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__147_i_7
       (.I0(alu_io_in1[12]),
        .I1(alu_io_in1[49]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [13]));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__148_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__148_i_4_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[51]_1 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__148_i_2
       (.I0(alu_io_in2[50]),
        .I1(alu_io_in1[50]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[51]_3 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__148_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_8),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[50]),
        .I4(alu_io_in2[50]),
        .I5(Q),
        .O(\bypass_mux_1_reg[51]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__148_i_4
       (.I0(core__145_i_7_n_0),
        .I1(core__147_i_5_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__146_i_5_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__148_i_5_n_0),
        .O(core__148_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__148_i_5
       (.I0(core__136_i_8_n_0),
        .I1(core__144_i_6_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__140_i_8_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__148_i_6_n_0),
        .O(core__148_i_5_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__148_i_6
       (.I0(core__641_i_12_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [44]),
        .I3(shamt),
        .I4(\alu/shin [12]),
        .O(core__148_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1800" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__148_i_7
       (.I0(alu_io_in1[11]),
        .I1(alu_io_in1[50]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [12]));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__149_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__149_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[52]_1 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__149_i_2
       (.I0(alu_io_in2[51]),
        .I1(alu_io_in1[51]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[52]_3 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__149_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_9),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[51]),
        .I4(alu_io_in2[51]),
        .I5(Q),
        .O(\bypass_mux_1_reg[52]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__149_i_5
       (.I0(core__146_i_5_n_0),
        .I1(core__148_i_5_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__147_i_5_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__149_i_6_n_0),
        .O(core__149_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__149_i_6
       (.I0(core__137_i_9_n_0),
        .I1(ex_ctrl_alu_dw_reg_33),
        .I2(alu_io_in2[2]),
        .I3(core__141_i_8_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__149_i_7_n_0),
        .O(core__149_i_6_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__149_i_7
       (.I0(core__639_i_10_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [43]),
        .I3(shamt),
        .I4(\alu/shin [11]),
        .O(core__149_i_7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1799" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__149_i_8
       (.I0(alu_io_in1[10]),
        .I1(alu_io_in1[51]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [11]));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__150_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__150_i_4_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[53]_1 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__150_i_2
       (.I0(alu_io_in2[52]),
        .I1(alu_io_in1[52]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[53]_3 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__150_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_10),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[52]),
        .I4(alu_io_in2[52]),
        .I5(Q),
        .O(\bypass_mux_1_reg[53]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__150_i_4
       (.I0(core__147_i_5_n_0),
        .I1(core__149_i_6_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__148_i_5_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__150_i_5_n_0),
        .O(core__150_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__150_i_5
       (.I0(core__138_i_8_n_0),
        .I1(core__146_i_6_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__142_i_7_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__150_i_6_n_0),
        .O(core__150_i_5_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__150_i_6
       (.I0(core__134_i_10_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [42]),
        .I3(shamt),
        .I4(\alu/shin [10]),
        .O(core__150_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1798" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__150_i_7
       (.I0(alu_io_in1[9]),
        .I1(alu_io_in1[52]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [10]));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__151_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__151_i_4_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[54]_1 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__151_i_2
       (.I0(alu_io_in2[53]),
        .I1(alu_io_in1[53]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[54]_3 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__151_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_11),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[53]),
        .I4(alu_io_in2[53]),
        .I5(Q),
        .O(\bypass_mux_1_reg[54]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__151_i_4
       (.I0(core__148_i_5_n_0),
        .I1(core__150_i_5_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__149_i_6_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__151_i_5_n_0),
        .O(core__151_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__151_i_5
       (.I0(core__139_i_8_n_0),
        .I1(core__147_i_6_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__143_i_7_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__151_i_6_n_0),
        .O(core__151_i_5_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__151_i_6
       (.I0(core__135_i_10_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [41]),
        .I3(shamt),
        .I4(\alu/shin [9]),
        .O(core__151_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1797" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__151_i_7
       (.I0(alu_io_in1[8]),
        .I1(alu_io_in1[53]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [9]));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__152_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__152_i_4_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[55]_1 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__152_i_2
       (.I0(alu_io_in2[54]),
        .I1(alu_io_in1[54]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[55]_3 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__152_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_12),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[54]),
        .I4(alu_io_in2[54]),
        .I5(Q),
        .O(\bypass_mux_1_reg[55]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__152_i_4
       (.I0(core__149_i_6_n_0),
        .I1(core__151_i_5_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__150_i_5_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__152_i_5_n_0),
        .O(core__152_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__152_i_5
       (.I0(core__140_i_8_n_0),
        .I1(core__148_i_6_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__144_i_6_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__152_i_6_n_0),
        .O(core__152_i_5_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__152_i_6
       (.I0(core__136_i_10_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [40]),
        .I3(shamt),
        .I4(\alu/shin [8]),
        .O(core__152_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1796" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__152_i_7
       (.I0(alu_io_in1[7]),
        .I1(alu_io_in1[54]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [8]));
  (* SOFT_HLUTNM = "soft_lutpair1814" *) 
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__153_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__153_i_5_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[56]_1 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__153_i_2
       (.I0(alu_io_in2[55]),
        .I1(alu_io_in1[55]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[56]_3 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__153_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_13),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[55]),
        .I4(alu_io_in2[55]),
        .I5(Q),
        .O(\bypass_mux_1_reg[56]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__153_i_5
       (.I0(core__150_i_5_n_0),
        .I1(core__152_i_5_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__151_i_5_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__153_i_6_n_0),
        .O(core__153_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__153_i_6
       (.I0(core__141_i_8_n_0),
        .I1(core__149_i_7_n_0),
        .I2(alu_io_in2[2]),
        .I3(ex_ctrl_alu_dw_reg_33),
        .I4(alu_io_in2[3]),
        .I5(core__153_i_7_n_0),
        .O(core__153_i_6_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__153_i_7
       (.I0(core__137_i_10_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [39]),
        .I3(shamt),
        .I4(\alu/shin [7]),
        .O(core__153_i_7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1795" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__153_i_8
       (.I0(alu_io_in1[6]),
        .I1(alu_io_in1[55]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [7]));
  LUT6 #(
    .INIT(64'hBBBFFFBFFFFFFFFF)) 
    core__154_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__154_i_4_n_0),
        .I3(alu_io_in2[0]),
        .I4(core__154_i_5_n_0),
        .I5(core__154_i_6_n_0),
        .O(\bypass_mux_1_reg[57]_1 ));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__154_i_10
       (.I0(\alu/shin [38]),
        .I1(shamt),
        .I2(alu_io_in1[5]),
        .I3(core__154_i_12_n_0),
        .I4(\alu/_T_55 ),
        .O(core__154_i_10_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1810" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__154_i_11
       (.I0(alu_io_in1[40]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__154_i_11_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1872" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__154_i_12
       (.I0(alu_io_in1[56]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__154_i_12_n_0));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__154_i_2
       (.I0(alu_io_in2[56]),
        .I1(alu_io_in1[56]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[57]_3 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__154_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_14),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[56]),
        .I4(alu_io_in2[56]),
        .I5(Q),
        .O(\bypass_mux_1_reg[57]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__154_i_4
       (.I0(core__152_i_5_n_0),
        .I1(alu_io_in2[1]),
        .I2(core__154_i_7_n_0),
        .I3(alu_io_in2[2]),
        .I4(core__154_i_8_n_0),
        .O(core__154_i_4_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1881" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__154_i_5
       (.I0(core__151_i_5_n_0),
        .I1(alu_io_in2[1]),
        .I2(core__153_i_6_n_0),
        .O(core__154_i_5_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1814" *) 
  LUT2 #(
    .INIT(4'h1)) 
    core__154_i_6
       (.I0(ex_ctrl_alu_fn[2]),
        .I1(Q),
        .O(core__154_i_6_n_0));
  LUT3 #(
    .INIT(8'hB8)) 
    core__154_i_7
       (.I0(core__142_i_7_n_0),
        .I1(alu_io_in2[3]),
        .I2(core__150_i_6_n_0),
        .O(core__154_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__154_i_8
       (.I0(core__146_i_6_n_0),
        .I1(alu_io_in2[3]),
        .I2(core__154_i_9_n_0),
        .I3(alu_io_in2[4]),
        .I4(core__154_i_10_n_0),
        .O(core__154_i_8_n_0));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__154_i_9
       (.I0(\alu/shin [54]),
        .I1(shamt),
        .I2(alu_io_in1[21]),
        .I3(core__154_i_11_n_0),
        .I4(\alu/_T_55 ),
        .O(core__154_i_9_n_0));
  LUT6 #(
    .INIT(64'hBBBFFFBFFFFFFFFF)) 
    core__155_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__155_i_4_n_0),
        .I3(alu_io_in2[0]),
        .I4(core__154_i_4_n_0),
        .I5(core__154_i_6_n_0),
        .O(\bypass_mux_1_reg[58]_1 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__155_i_2
       (.I0(alu_io_in2[57]),
        .I1(alu_io_in1[57]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[58]_3 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__155_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_15),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[57]),
        .I4(alu_io_in2[57]),
        .I5(Q),
        .O(\bypass_mux_1_reg[58]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1881" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__155_i_4
       (.I0(core__153_i_6_n_0),
        .I1(alu_io_in2[1]),
        .I2(core__155_i_5_n_0),
        .O(core__155_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__155_i_5
       (.I0(core__143_i_7_n_0),
        .I1(core__151_i_6_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__147_i_6_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__155_i_6_n_0),
        .O(core__155_i_5_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__155_i_6
       (.I0(core__159_i_8_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [37]),
        .I3(shamt),
        .I4(\alu/shin [5]),
        .O(core__155_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1793" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__155_i_7
       (.I0(alu_io_in1[4]),
        .I1(alu_io_in1[57]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [5]));
  LUT6 #(
    .INIT(64'hBBBFFFBFFFFFFFFF)) 
    core__156_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__156_i_4_n_0),
        .I3(alu_io_in2[0]),
        .I4(core__155_i_4_n_0),
        .I5(core__154_i_6_n_0),
        .O(\bypass_mux_1_reg[59]_1 ));
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    core__156_i_2
       (.I0(alu_io_in2[58]),
        .I1(alu_io_in1[58]),
        .I2(Q),
        .I3(ex_ctrl_alu_fn[2]),
        .I4(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[59]_3 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__156_i_3
       (.I0(\alu/_T_55 ),
        .I1(ex_reg_rvc_reg_16),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[58]),
        .I4(alu_io_in2[58]),
        .I5(Q),
        .O(\bypass_mux_1_reg[59]_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__156_i_4
       (.I0(core__154_i_7_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__154_i_8_n_0),
        .I3(alu_io_in2[1]),
        .I4(core__156_i_5_n_0),
        .O(core__156_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__156_i_5
       (.I0(core__144_i_6_n_0),
        .I1(core__152_i_6_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__148_i_6_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__156_i_6_n_0),
        .O(core__156_i_5_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__156_i_6
       (.I0(core__140_i_9_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [36]),
        .I3(shamt),
        .I4(\alu/shin [4]),
        .O(core__156_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1792" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__156_i_7
       (.I0(alu_io_in1[3]),
        .I1(alu_io_in1[58]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [4]));
  LUT6 #(
    .INIT(64'hBBBFFFBFFFFFFFFF)) 
    core__157_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__157_i_4_n_0),
        .I3(alu_io_in2[0]),
        .I4(core__156_i_4_n_0),
        .I5(core__154_i_6_n_0),
        .O(\bypass_mux_1_reg[60]_1 ));
  LUT6 #(
    .INIT(64'h1CC35FFF00000000)) 
    core__157_i_2
       (.I0(\alu/_T_205 ),
        .I1(Q),
        .I2(alu_io_in2[59]),
        .I3(alu_io_in1[59]),
        .I4(\alu/_T_198 ),
        .I5(core__157_i_5_n_0),
        .O(\bypass_mux_1_reg[60]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1880" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__157_i_4
       (.I0(core__155_i_5_n_0),
        .I1(alu_io_in2[1]),
        .I2(core__157_i_6_n_0),
        .O(core__157_i_4_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1885" *) 
  LUT2 #(
    .INIT(4'h7)) 
    core__157_i_5
       (.I0(\ex_ctrl_alu_fn_reg[3]_6 ),
        .I1(\alu/_T_55 ),
        .O(core__157_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__157_i_6
       (.I0(ex_ctrl_alu_dw_reg_33),
        .I1(core__153_i_7_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__149_i_7_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__157_i_7_n_0),
        .O(core__157_i_6_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__157_i_7
       (.I0(core__141_i_9_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [35]),
        .I3(shamt),
        .I4(\alu/shin [3]),
        .O(core__157_i_7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1788" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__157_i_8
       (.I0(alu_io_in1[2]),
        .I1(alu_io_in1[59]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [3]));
  (* SOFT_HLUTNM = "soft_lutpair1802" *) 
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__158_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__158_i_3_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(\bypass_mux_1_reg[61]_1 ));
  LUT6 #(
    .INIT(64'h1CC35FFF00000000)) 
    core__158_i_2
       (.I0(\alu/_T_205 ),
        .I1(Q),
        .I2(alu_io_in2[60]),
        .I3(alu_io_in1[60]),
        .I4(\alu/_T_198 ),
        .I5(core__158_i_4_n_0),
        .O(\bypass_mux_1_reg[61]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__158_i_3
       (.I0(core__155_i_5_n_0),
        .I1(core__157_i_6_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__156_i_5_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__158_i_5_n_0),
        .O(core__158_i_3_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    core__158_i_4
       (.I0(\ex_ctrl_alu_fn_reg[3]_7 ),
        .I1(\alu/_T_55 ),
        .O(core__158_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__158_i_5
       (.I0(core__146_i_6_n_0),
        .I1(core__158_i_6_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__150_i_6_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__158_i_7_n_0),
        .O(core__158_i_5_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__158_i_6
       (.I0(core__154_i_9_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [38]),
        .I3(shamt),
        .I4(\alu/shin [6]),
        .O(core__158_i_6_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__158_i_7
       (.I0(core__142_i_8_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [34]),
        .I3(shamt),
        .I4(\alu/shin [2]),
        .O(core__158_i_7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1794" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__158_i_8
       (.I0(alu_io_in1[5]),
        .I1(alu_io_in1[56]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [6]));
  (* SOFT_HLUTNM = "soft_lutpair1784" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__158_i_9
       (.I0(alu_io_in1[1]),
        .I1(alu_io_in1[60]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [2]));
  LUT6 #(
    .INIT(64'hBBBFFFBFFFFFFFFF)) 
    core__159_i_1
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__159_i_3_n_0),
        .I3(alu_io_in2[0]),
        .I4(core__159_i_4_n_0),
        .I5(core__154_i_6_n_0),
        .O(\bypass_mux_1_reg[62]_1 ));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__159_i_10
       (.I0(\alu/shin [49]),
        .I1(shamt),
        .I2(alu_io_in1[16]),
        .I3(core__159_i_14_n_0),
        .I4(\alu/_T_55 ),
        .O(core__159_i_10_n_0));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__159_i_11
       (.I0(\alu/shin [33]),
        .I1(shamt),
        .I2(alu_io_in1[0]),
        .I3(core__159_i_15_n_0),
        .I4(\alu/_T_55 ),
        .O(core__159_i_11_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1811" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__159_i_12
       (.I0(alu_io_in1[41]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__159_i_12_n_0));
  LUT3 #(
    .INIT(8'hB8)) 
    core__159_i_13
       (.I0(alu_io_in1[57]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__159_i_13_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1806" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__159_i_14
       (.I0(alu_io_in1[45]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__159_i_14_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1872" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__159_i_15
       (.I0(alu_io_in1[61]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__159_i_15_n_0));
  LUT6 #(
    .INIT(64'h1CC35FFF00000000)) 
    core__159_i_2
       (.I0(\alu/_T_205 ),
        .I1(Q),
        .I2(alu_io_in2[61]),
        .I3(alu_io_in1[61]),
        .I4(\alu/_T_198 ),
        .I5(core__159_i_5_n_0),
        .O(\bypass_mux_1_reg[62]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__159_i_3
       (.I0(core__157_i_6_n_0),
        .I1(alu_io_in2[1]),
        .I2(core__159_i_6_n_0),
        .I3(alu_io_in2[2]),
        .I4(core__159_i_7_n_0),
        .O(core__159_i_3_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1880" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__159_i_4
       (.I0(core__156_i_5_n_0),
        .I1(alu_io_in2[1]),
        .I2(core__158_i_5_n_0),
        .O(core__159_i_4_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1885" *) 
  LUT2 #(
    .INIT(4'h7)) 
    core__159_i_5
       (.I0(\bypass_mux_1[1]_i_5_n_0 ),
        .I1(\alu/_T_55 ),
        .O(core__159_i_5_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__159_i_6
       (.I0(core__147_i_6_n_0),
        .I1(alu_io_in2[3]),
        .I2(core__159_i_8_n_0),
        .I3(alu_io_in2[4]),
        .I4(core__159_i_9_n_0),
        .O(core__159_i_6_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__159_i_7
       (.I0(core__151_i_6_n_0),
        .I1(alu_io_in2[3]),
        .I2(core__159_i_10_n_0),
        .I3(alu_io_in2[4]),
        .I4(core__159_i_11_n_0),
        .O(core__159_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__159_i_8
       (.I0(\alu/shin [53]),
        .I1(shamt),
        .I2(alu_io_in1[20]),
        .I3(core__159_i_12_n_0),
        .I4(\alu/_T_55 ),
        .O(core__159_i_8_n_0));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__159_i_9
       (.I0(\alu/shin [37]),
        .I1(shamt),
        .I2(alu_io_in1[4]),
        .I3(core__159_i_13_n_0),
        .I4(\alu/_T_55 ),
        .O(core__159_i_9_n_0));
  LUT6 #(
    .INIT(64'h5555555557555555)) 
    core__160_i_1
       (.I0(core__160_i_2_n_0),
        .I1(ex_ctrl_alu_fn[2]),
        .I2(Q),
        .I3(core__160_i_3_n_0),
        .I4(ex_ctrl_alu_fn[0]),
        .I5(ex_ctrl_alu_fn[1]),
        .O(\bypass_mux_1_reg[63]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1840" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__160_i_10
       (.I0(\bypass_mux_1_reg[0]_0 ),
        .I1(alu_io_in1[62]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [0]));
  LUT6 #(
    .INIT(64'h1CC35FFF00000000)) 
    core__160_i_2
       (.I0(\alu/_T_205 ),
        .I1(Q),
        .I2(alu_io_in2[62]),
        .I3(alu_io_in1[62]),
        .I4(\alu/_T_198 ),
        .I5(core__160_i_4_n_0),
        .O(core__160_i_2_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__160_i_3
       (.I0(core__157_i_6_n_0),
        .I1(core__160_i_5_n_0),
        .I2(alu_io_in2[0]),
        .I3(core__158_i_5_n_0),
        .I4(alu_io_in2[1]),
        .I5(core__160_i_6_n_0),
        .O(core__160_i_3_n_0));
  LUT5 #(
    .INIT(32'h0F1DFFFF)) 
    core__160_i_4
       (.I0(\bypass_mux_1_reg[1]_1 ),
        .I1(alu_io_in2[1]),
        .I2(_T_121),
        .I3(alu_io_in2[0]),
        .I4(\alu/_T_55 ),
        .O(core__160_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__160_i_5
       (.I0(core__147_i_6_n_0),
        .I1(core__155_i_6_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__151_i_6_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__160_i_7_n_0),
        .O(core__160_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__160_i_6
       (.I0(core__148_i_6_n_0),
        .I1(core__156_i_6_n_0),
        .I2(alu_io_in2[2]),
        .I3(core__152_i_6_n_0),
        .I4(alu_io_in2[3]),
        .I5(core__160_i_8_n_0),
        .O(core__160_i_6_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__160_i_7
       (.I0(core__159_i_10_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [33]),
        .I3(shamt),
        .I4(\alu/shin [1]),
        .O(core__160_i_7_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    core__160_i_8
       (.I0(core__144_i_7_n_0),
        .I1(alu_io_in2[4]),
        .I2(\alu/shin [32]),
        .I3(shamt),
        .I4(\alu/shin [0]),
        .O(core__160_i_8_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1791" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__160_i_9
       (.I0(alu_io_in1[0]),
        .I1(alu_io_in1[61]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [1]));
  LUT5 #(
    .INIT(32'hEAAAFFFF)) 
    core__161_i_2
       (.I0(core__161_i_3_n_0),
        .I1(alu_io_in2[30]),
        .I2(alu_io_in1[30]),
        .I3(\alu/_T_205 ),
        .I4(core__161_i_4_n_0),
        .O(\bypass_mux_1_reg[32]_0 ));
  LUT6 #(
    .INIT(64'hF88888F888F8F888)) 
    core__161_i_3
       (.I0(\alu/_T_55 ),
        .I1(core__161_i_5_n_0),
        .I2(\alu/_T_198 ),
        .I3(alu_io_in1[30]),
        .I4(alu_io_in2[30]),
        .I5(Q),
        .O(core__161_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    core__161_i_4
       (.I0(ex_ctrl_alu_fn[1]),
        .I1(ex_ctrl_alu_fn[0]),
        .I2(core__161_i_6_n_0),
        .I3(Q),
        .I4(ex_ctrl_alu_fn[2]),
        .O(core__161_i_4_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__161_i_5
       (.I0(\bypass_mux_1_reg[29]_0 ),
        .I1(\bypass_mux_1_reg[34]_2 ),
        .I2(alu_io_in2[0]),
        .I3(\bypass_mux_1_reg[33]_2 ),
        .I4(alu_io_in2[1]),
        .I5(\bypass_mux_1_reg[35]_2 ),
        .O(core__161_i_5_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__161_i_6
       (.I0(\bypass_mux_1_reg[29]_1 ),
        .I1(\bypass_mux_1_reg[33]_2 ),
        .I2(alu_io_in2[0]),
        .I3(\bypass_mux_1_reg[29]_0 ),
        .I4(alu_io_in2[1]),
        .I5(\bypass_mux_1_reg[34]_2 ),
        .O(core__161_i_6_n_0));
  LUT4 #(
    .INIT(16'h3808)) 
    core__162_i_1
       (.I0(div_n_138),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[1]),
        .O(alu_io_in1[0]));
  LUT5 #(
    .INIT(32'hCFECCCEC)) 
    core__162_i_2
       (.I0(mem_reg_rvc_reg_0),
        .I1(core__162_i_5_n_0),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(ex_ctrl_sel_alu2[1]),
        .I4(\divisor_reg[57] [0]),
        .O(alu_io_in2[1]));
  LUT4 #(
    .INIT(16'h30A0)) 
    core__162_i_3
       (.I0(mem_reg_rs2[0]),
        .I1(core__162_i_6_n_0),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(ex_ctrl_sel_alu2[0]),
        .O(alu_io_in2[0]));
  (* SOFT_HLUTNM = "soft_lutpair1857" *) 
  LUT3 #(
    .INIT(8'h08)) 
    core__162_i_4
       (.I0(div_n_240),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .O(\bypass_mux_1_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFF00B8000000B800)) 
    core__162_i_5
       (.I0(\ex_reg_inst_reg_n_0_[16] ),
        .I1(\ex_ctrl_sel_imm_reg[1]_1 ),
        .I2(\ex_reg_inst_reg_n_0_[21] ),
        .I3(core__163_i_6_n_0),
        .I4(core__163_i_5_n_0),
        .I5(\mem_reg_inst_reg[31]_0 [1]),
        .O(core__162_i_5_n_0));
  LUT6 #(
    .INIT(64'hFFFF55FFFFFF330F)) 
    core__162_i_6
       (.I0(\ex_reg_inst_reg_n_0_[15] ),
        .I1(_T_1710),
        .I2(\mem_reg_inst_reg[31]_0 [0]),
        .I3(\bypass_mux_1_reg[6]_1 [2]),
        .I4(\bypass_mux_1_reg[6]_1 [1]),
        .I5(\bypass_mux_1_reg[6]_1 [0]),
        .O(core__162_i_6_n_0));
  LUT4 #(
    .INIT(16'h3808)) 
    core__163_i_1
       (.I0(div_n_141),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[4]),
        .O(alu_io_in1[3]));
  LUT6 #(
    .INIT(64'hF4FF444444444444)) 
    core__163_i_2
       (.I0(\bypass_mux_1_reg[4]_0 ),
        .I1(mem_reg_rs2[4]),
        .I2(\mem_reg_inst_reg[31]_0 [4]),
        .I3(core__163_i_5_n_0),
        .I4(core__163_i_6_n_0),
        .I5(core__163_i_7_n_0),
        .O(alu_io_in2[4]));
  LUT6 #(
    .INIT(64'hF4FF444444444444)) 
    core__163_i_3
       (.I0(\bypass_mux_1_reg[4]_0 ),
        .I1(mem_reg_rs2[3]),
        .I2(\mem_reg_inst_reg[31]_0 [3]),
        .I3(core__163_i_5_n_0),
        .I4(core__163_i_6_n_0),
        .I5(core__163_i_8_n_0),
        .O(alu_io_in2[3]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__163_i_4
       (.I0(div_n_140),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[3]),
        .O(alu_io_in1[2]));
  (* SOFT_HLUTNM = "soft_lutpair1822" *) 
  LUT2 #(
    .INIT(4'h1)) 
    core__163_i_5
       (.I0(\bypass_mux_1_reg[6]_1 [1]),
        .I1(\bypass_mux_1_reg[6]_1 [2]),
        .O(core__163_i_5_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1790" *) 
  LUT5 #(
    .INIT(32'h88888088)) 
    core__163_i_6
       (.I0(ex_ctrl_sel_alu2[0]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(\bypass_mux_1_reg[6]_1 [0]),
        .I3(\bypass_mux_1_reg[6]_1 [1]),
        .I4(\bypass_mux_1_reg[6]_1 [2]),
        .O(core__163_i_6_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1822" *) 
  LUT5 #(
    .INIT(32'hAAEFAA2F)) 
    core__163_i_7
       (.I0(\ex_reg_inst_reg_n_0_[24] ),
        .I1(\bypass_mux_1_reg[6]_1 [0]),
        .I2(\bypass_mux_1_reg[6]_1 [2]),
        .I3(\bypass_mux_1_reg[6]_1 [1]),
        .I4(\ex_reg_inst_reg_n_0_[19] ),
        .O(core__163_i_7_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1787" *) 
  LUT5 #(
    .INIT(32'hAAEFAA2F)) 
    core__163_i_8
       (.I0(\ex_reg_inst_reg_n_0_[23] ),
        .I1(\bypass_mux_1_reg[6]_1 [0]),
        .I2(\bypass_mux_1_reg[6]_1 [2]),
        .I3(\bypass_mux_1_reg[6]_1 [1]),
        .I4(\ex_reg_inst_reg_n_0_[18] ),
        .O(core__163_i_8_n_0));
  LUT4 #(
    .INIT(16'h3808)) 
    core__164_i_1
       (.I0(div_n_145),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[8]),
        .O(alu_io_in1[7]));
  LUT5 #(
    .INIT(32'h04FF0404)) 
    core__164_i_2
       (.I0(ex_ctrl_sel_alu2[0]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(div_n_218),
        .I3(\bypass_mux_1_reg[6]_0 ),
        .I4(\ex_reg_inst_reg_n_0_[28] ),
        .O(alu_io_in2[7]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__164_i_3
       (.I0(div_n_144),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[7]),
        .O(alu_io_in1[6]));
  LUT5 #(
    .INIT(32'h40FF4040)) 
    core__164_i_4
       (.I0(ex_ctrl_sel_alu2[0]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(\divisor_reg[57] [2]),
        .I3(\bypass_mux_1_reg[6]_0 ),
        .I4(\mem_reg_inst_reg[31]_0 [6]),
        .O(alu_io_in2[6]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__165_i_1
       (.I0(div_n_147),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[10]),
        .O(alu_io_in1[9]));
  LUT5 #(
    .INIT(32'h04FF0404)) 
    core__165_i_2
       (.I0(ex_ctrl_sel_alu2[0]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(div_n_219),
        .I3(\bypass_mux_1_reg[6]_0 ),
        .I4(\ex_reg_inst_reg_n_0_[30] ),
        .O(alu_io_in2[9]));
  LUT5 #(
    .INIT(32'h04FF0404)) 
    core__165_i_3
       (.I0(ex_ctrl_sel_alu2[0]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(\mem_reg_rs2_reg[25]_0 ),
        .I3(\bypass_mux_1_reg[6]_0 ),
        .I4(\ex_reg_inst_reg_n_0_[29] ),
        .O(alu_io_in2[8]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__165_i_4
       (.I0(div_n_146),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[9]),
        .O(alu_io_in1[8]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__166_i_1
       (.I0(div_n_151),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[14]),
        .O(alu_io_in1[13]));
  LUT6 #(
    .INIT(64'hC404C4C4C4040404)) 
    core__166_i_2
       (.I0(div_n_223),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[14] ),
        .I4(core__166_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[13]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__166_i_3
       (.I0(div_n_150),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[13]),
        .O(alu_io_in1[12]));
  LUT6 #(
    .INIT(64'hC404C4C4C4040404)) 
    core__166_i_4
       (.I0(div_n_222),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[13] ),
        .I4(core__166_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[12]));
  (* SOFT_HLUTNM = "soft_lutpair1846" *) 
  LUT2 #(
    .INIT(4'h2)) 
    core__166_i_5
       (.I0(\bypass_mux_1_reg[6]_1 [1]),
        .I1(\bypass_mux_1_reg[6]_1 [2]),
        .O(core__166_i_5_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1846" *) 
  LUT4 #(
    .INIT(16'hAA2A)) 
    core__166_i_6
       (.I0(\mem_reg_inst_reg[31]_0 [7]),
        .I1(\bypass_mux_1_reg[6]_1 [0]),
        .I2(\bypass_mux_1_reg[6]_1 [2]),
        .I3(\bypass_mux_1_reg[6]_1 [1]),
        .O(core__166_i_6_n_0));
  LUT4 #(
    .INIT(16'h3808)) 
    core__167_i_1
       (.I0(div_n_154),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[17]),
        .O(alu_io_in1[16]));
  LUT6 #(
    .INIT(64'hC808C8C8C8080808)) 
    core__167_i_2
       (.I0(mem_reg_rs2[17]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[17] ),
        .I4(core__166_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[16]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__167_i_3
       (.I0(div_n_153),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[16]),
        .O(alu_io_in1[15]));
  LUT6 #(
    .INIT(64'hC808C8C8C8080808)) 
    core__167_i_4
       (.I0(mem_reg_rs2[16]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[16] ),
        .I4(core__166_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[15]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__168_i_1
       (.I0(div_n_157),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[20]),
        .O(alu_io_in1[19]));
  LUT6 #(
    .INIT(64'hC404C4C4C4040404)) 
    core__168_i_2
       (.I0(div_n_227),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(_T_1710),
        .I4(core__168_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[19]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__168_i_3
       (.I0(div_n_156),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[19]),
        .O(alu_io_in1[18]));
  LUT6 #(
    .INIT(64'hC404C4C4C4040404)) 
    core__168_i_4
       (.I0(div_n_226),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[19] ),
        .I4(core__166_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[18]));
  (* SOFT_HLUTNM = "soft_lutpair1787" *) 
  LUT3 #(
    .INIT(8'h04)) 
    core__168_i_5
       (.I0(\bypass_mux_1_reg[6]_1 [2]),
        .I1(\bypass_mux_1_reg[6]_1 [1]),
        .I2(\bypass_mux_1_reg[6]_1 [0]),
        .O(core__168_i_5_n_0));
  LUT4 #(
    .INIT(16'h3808)) 
    core__169_i_1
       (.I0(div_n_160),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[23]),
        .O(alu_io_in1[22]));
  LUT6 #(
    .INIT(64'hC404C4C4C4040404)) 
    core__169_i_2
       (.I0(div_n_230),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[23] ),
        .I4(core__168_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[22]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__169_i_3
       (.I0(div_n_159),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[22]),
        .O(alu_io_in1[21]));
  LUT6 #(
    .INIT(64'hC404C4C4C4040404)) 
    core__169_i_4
       (.I0(div_n_229),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[22] ),
        .I4(core__168_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[21]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__170_i_1
       (.I0(div_n_163),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[26]),
        .O(alu_io_in1[25]));
  LUT6 #(
    .INIT(64'hC808C8C8C8080808)) 
    core__170_i_2
       (.I0(mem_reg_rs2[26]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\mem_reg_inst_reg[31]_0 [5]),
        .I4(core__168_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[25]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__170_i_3
       (.I0(div_n_162),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[25]),
        .O(alu_io_in1[24]));
  LUT6 #(
    .INIT(64'hC808C8C8C8080808)) 
    core__170_i_4
       (.I0(\divisor_reg[57] [3]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[25] ),
        .I4(core__168_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[24]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__171_i_1
       (.I0(div_n_166),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[29]),
        .O(alu_io_in1[28]));
  LUT6 #(
    .INIT(64'hC808C8C8C8080808)) 
    core__171_i_2
       (.I0(mem_reg_rs2[29]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[29] ),
        .I4(core__168_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[28]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__171_i_3
       (.I0(div_n_165),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[28]),
        .O(alu_io_in1[27]));
  LUT6 #(
    .INIT(64'hC808C8C8C8080808)) 
    core__171_i_4
       (.I0(mem_reg_rs2[28]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[28] ),
        .I4(core__168_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[27]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__172_i_1
       (.I0(div_n_170),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[32]),
        .O(alu_io_in1[31]));
  (* SOFT_HLUTNM = "soft_lutpair1844" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__172_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[32]),
        .O(alu_io_in2[31]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__172_i_3
       (.I0(\remainder_reg[31] ),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(\mem_reg_pc_reg[31]_0 ),
        .O(alu_io_in1[30]));
  (* SOFT_HLUTNM = "soft_lutpair1858" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__172_i_4
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[31]),
        .O(alu_io_in2[30]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__173_i_1
       (.I0(\remainder_reg[35]_0 ),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[35]),
        .O(alu_io_in1[34]));
  (* SOFT_HLUTNM = "soft_lutpair1848" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__173_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[35]),
        .O(alu_io_in2[34]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__173_i_3
       (.I0(\remainder_reg[34]_0 ),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[34]),
        .O(alu_io_in1[33]));
  (* SOFT_HLUTNM = "soft_lutpair1850" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__173_i_4
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[34]),
        .O(alu_io_in2[33]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__174_i_1
       (.I0(\remainder_reg[38]_0 ),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[38]),
        .O(alu_io_in1[37]));
  (* SOFT_HLUTNM = "soft_lutpair1853" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__174_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[38]),
        .O(alu_io_in2[37]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__174_i_3
       (.I0(\remainder_reg[37]_0 ),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[37]),
        .O(alu_io_in1[36]));
  (* SOFT_HLUTNM = "soft_lutpair1845" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__174_i_4
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[37]),
        .O(alu_io_in2[36]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__175_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [1]),
        .O(alu_io_in1[40]));
  (* SOFT_HLUTNM = "soft_lutpair1844" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__175_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(\divisor_reg[57] [4]),
        .O(alu_io_in2[40]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__175_i_3
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(_T_2770[1]),
        .O(alu_io_in1[39]));
  (* SOFT_HLUTNM = "soft_lutpair1851" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__175_i_4
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[40]),
        .O(alu_io_in2[39]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__176_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [4]),
        .O(alu_io_in1[43]));
  (* SOFT_HLUTNM = "soft_lutpair1855" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__176_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[44]),
        .O(alu_io_in2[43]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__176_i_3
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [3]),
        .O(alu_io_in1[42]));
  (* SOFT_HLUTNM = "soft_lutpair1856" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__176_i_4
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[43]),
        .O(alu_io_in2[42]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__177_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [6]),
        .O(alu_io_in1[46]));
  (* SOFT_HLUTNM = "soft_lutpair1852" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__177_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[47]),
        .O(alu_io_in2[46]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__177_i_3
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [5]),
        .O(alu_io_in1[45]));
  (* SOFT_HLUTNM = "soft_lutpair1859" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__177_i_4
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[46]),
        .O(alu_io_in2[45]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__178_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [8]),
        .O(alu_io_in1[49]));
  (* SOFT_HLUTNM = "soft_lutpair1856" *) 
  LUT4 #(
    .INIT(16'hAABA)) 
    core__178_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(div_n_234),
        .O(alu_io_in2[49]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__178_i_3
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [7]),
        .O(alu_io_in1[48]));
  (* SOFT_HLUTNM = "soft_lutpair1847" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__178_i_4
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[49]),
        .O(alu_io_in2[48]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__179_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(_T_2770[14]),
        .O(alu_io_in1[52]));
  (* SOFT_HLUTNM = "soft_lutpair1853" *) 
  LUT4 #(
    .INIT(16'hAABA)) 
    core__179_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(div_n_237),
        .O(alu_io_in2[52]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__179_i_3
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [10]),
        .O(alu_io_in1[51]));
  (* SOFT_HLUTNM = "soft_lutpair1854" *) 
  LUT4 #(
    .INIT(16'hAABA)) 
    core__179_i_4
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(div_n_236),
        .O(alu_io_in2[51]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__180_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(_T_2770[17]),
        .O(alu_io_in1[55]));
  (* SOFT_HLUTNM = "soft_lutpair1860" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__180_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[56]),
        .O(alu_io_in2[55]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__180_i_3
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [12]),
        .O(alu_io_in1[54]));
  (* SOFT_HLUTNM = "soft_lutpair1860" *) 
  LUT4 #(
    .INIT(16'hAABA)) 
    core__180_i_4
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(div_n_239),
        .O(alu_io_in2[54]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__181_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(_T_2770[20]),
        .O(alu_io_in1[58]));
  (* SOFT_HLUTNM = "soft_lutpair1861" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__181_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[59]),
        .O(alu_io_in2[58]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__181_i_3
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [14]),
        .O(alu_io_in1[57]));
  (* SOFT_HLUTNM = "soft_lutpair1848" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__181_i_4
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[58]),
        .O(alu_io_in2[57]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__182_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [17]),
        .O(alu_io_in1[61]));
  (* SOFT_HLUTNM = "soft_lutpair1851" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__182_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[62]),
        .O(alu_io_in2[61]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__182_i_3
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [16]),
        .O(alu_io_in1[60]));
  (* SOFT_HLUTNM = "soft_lutpair1845" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__182_i_4
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[61]),
        .O(alu_io_in2[60]));
  LUT6 #(
    .INIT(64'h0000040000000000)) 
    core__193_i_1
       (.I0(\s1_req_cmd_reg[4] [0]),
        .I1(\s1_req_cmd_reg[4] [2]),
        .I2(\s1_req_cmd_reg[4] [1]),
        .I3(\s1_req_cmd_reg[4] [4]),
        .I4(\s1_req_cmd_reg[4] [3]),
        .I5(ex_ctrl_mem),
        .O(ex_sfence));
  (* SOFT_HLUTNM = "soft_lutpair1867" *) 
  LUT3 #(
    .INIT(8'h01)) 
    core__193_i_2
       (.I0(ex_reg_replay),
        .I1(ex_reg_valid),
        .I2(ex_reg_xcpt_interrupt),
        .O(mem_reg_sfence_reg_0));
  LUT5 #(
    .INIT(32'h00400000)) 
    core__196_i_1
       (.I0(\s1_req_cmd_reg[4] [3]),
        .I1(\s1_req_cmd_reg[4] [0]),
        .I2(\s1_req_cmd_reg[4] [2]),
        .I3(\s1_req_cmd_reg[4] [4]),
        .I4(\s1_req_cmd_reg[4] [1]),
        .O(mem_reg_slow_bypass_reg_0));
  (* SOFT_HLUTNM = "soft_lutpair1789" *) 
  LUT5 #(
    .INIT(32'hAAA20008)) 
    core__200_i_1
       (.I0(mem_ctrl_branch),
        .I1(\trig_state_reg[1]_1 ),
        .I2(\trig_state_reg[0]_0 ),
        .I3(\trig_state_reg[1]_0 ),
        .I4(mem_br_taken_),
        .O(\bypass_mux_2_reg[35]_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    core__266_i_10
       (.I0(\trig_pc_reg[63]_0 [49]),
        .I1(\trig_pc_reg[63]_0 [48]),
        .I2(\trig_pc_reg[63]_0 [50]),
        .O(\trig_pc_reg[0]_6 [0]));
  LUT3 #(
    .INIT(8'h01)) 
    core__266_i_12
       (.I0(\trig_pc_reg[63]_0 [46]),
        .I1(\trig_pc_reg[63]_0 [45]),
        .I2(\trig_pc_reg[63]_0 [47]),
        .O(\trig_pc_reg[0]_5 [3]));
  LUT3 #(
    .INIT(8'h01)) 
    core__266_i_13
       (.I0(\trig_pc_reg[63]_0 [43]),
        .I1(\trig_pc_reg[63]_0 [42]),
        .I2(\trig_pc_reg[63]_0 [44]),
        .O(\trig_pc_reg[0]_5 [2]));
  LUT4 #(
    .INIT(16'h1001)) 
    core__266_i_14
       (.I0(\trig_pc_reg[63]_0 [41]),
        .I1(\trig_pc_reg[63]_0 [40]),
        .I2(\trig_pc_reg[63]_0 [39]),
        .I3(\wb_reg_pc_reg[39]_0 [32]),
        .O(\trig_pc_reg[0]_5 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_15
       (.I0(\trig_pc_reg[63]_0 [38]),
        .I1(\wb_reg_pc_reg[39]_0 [31]),
        .I2(\wb_reg_pc_reg[39]_0 [29]),
        .I3(\trig_pc_reg[63]_0 [36]),
        .I4(\wb_reg_pc_reg[39]_0 [30]),
        .I5(\trig_pc_reg[63]_0 [37]),
        .O(\trig_pc_reg[0]_5 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_17
       (.I0(\trig_pc_reg[63]_0 [35]),
        .I1(\wb_reg_pc_reg[39]_0 [28]),
        .I2(\wb_reg_pc_reg[34]_0 [2]),
        .I3(\trig_pc_reg[63]_0 [33]),
        .I4(\wb_reg_pc_reg[34]_0 [3]),
        .I5(\trig_pc_reg[63]_0 [34]),
        .O(\trig_pc_reg[0]_4 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_18
       (.I0(\wb_reg_pc_reg[34]_0 [1]),
        .I1(\trig_pc_reg[63]_0 [32]),
        .I2(\bypass_mux_2_reg[31]_0 [2]),
        .I3(\trig_pc_reg[63]_0 [30]),
        .I4(\trig_pc_reg[63]_0 [31]),
        .I5(\wb_reg_pc_reg[39]_0 [27]),
        .O(\trig_pc_reg[0]_4 [2]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_19
       (.I0(\wb_reg_pc_reg[39]_0 [26]),
        .I1(\trig_pc_reg[63]_0 [27]),
        .I2(\bypass_mux_2_reg[31]_0 [0]),
        .I3(\trig_pc_reg[63]_0 [28]),
        .I4(\trig_pc_reg[63]_0 [29]),
        .I5(\bypass_mux_2_reg[31]_0 [1]),
        .O(\trig_pc_reg[0]_4 [1]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    core__266_i_2
       (.I0(mem_ctrl_jalr),
        .I1(trig_jalr_count_reg__0[2]),
        .I2(trig_jalr_count_reg__0[0]),
        .I3(trig_jalr_count_reg__0[1]),
        .I4(trig_jalr_count_reg__0[3]),
        .I5(trig_jalr_count_reg__0[4]),
        .O(\trig_pc_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_20
       (.I0(\wb_reg_pc_reg[39]_0 [23]),
        .I1(\trig_pc_reg[63]_0 [24]),
        .I2(\wb_reg_pc_reg[39]_0 [24]),
        .I3(\trig_pc_reg[63]_0 [25]),
        .I4(\trig_pc_reg[63]_0 [26]),
        .I5(\wb_reg_pc_reg[39]_0 [25]),
        .O(\trig_pc_reg[0]_4 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_22
       (.I0(\wb_reg_pc_reg[39]_0 [20]),
        .I1(\trig_pc_reg[63]_0 [21]),
        .I2(\wb_reg_pc_reg[39]_0 [21]),
        .I3(\trig_pc_reg[63]_0 [22]),
        .I4(\trig_pc_reg[63]_0 [23]),
        .I5(\wb_reg_pc_reg[39]_0 [22]),
        .O(\trig_pc_reg[0]_3 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_23
       (.I0(\wb_reg_pc_reg[39]_0 [17]),
        .I1(\trig_pc_reg[63]_0 [18]),
        .I2(\wb_reg_pc_reg[39]_0 [18]),
        .I3(\trig_pc_reg[63]_0 [19]),
        .I4(\trig_pc_reg[63]_0 [20]),
        .I5(\wb_reg_pc_reg[39]_0 [19]),
        .O(\trig_pc_reg[0]_3 [2]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_24
       (.I0(\wb_reg_pc_reg[39]_0 [16]),
        .I1(\trig_pc_reg[63]_0 [17]),
        .I2(\wb_reg_pc_reg[39]_0 [14]),
        .I3(\trig_pc_reg[63]_0 [15]),
        .I4(\trig_pc_reg[63]_0 [16]),
        .I5(\wb_reg_pc_reg[39]_0 [15]),
        .O(\trig_pc_reg[0]_3 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_25
       (.I0(\wb_reg_pc_reg[39]_0 [13]),
        .I1(\trig_pc_reg[63]_0 [14]),
        .I2(\wb_reg_pc_reg[39]_0 [11]),
        .I3(\trig_pc_reg[63]_0 [12]),
        .I4(\trig_pc_reg[63]_0 [13]),
        .I5(\wb_reg_pc_reg[39]_0 [12]),
        .O(\trig_pc_reg[0]_3 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_26
       (.I0(\wb_reg_pc_reg[39]_0 [8]),
        .I1(\trig_pc_reg[63]_0 [9]),
        .I2(\wb_reg_pc_reg[39]_0 [9]),
        .I3(\trig_pc_reg[63]_0 [10]),
        .I4(\trig_pc_reg[63]_0 [11]),
        .I5(\wb_reg_pc_reg[39]_0 [10]),
        .O(\trig_pc_reg[0]_2 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_27
       (.I0(\wb_reg_pc_reg[39]_0 [5]),
        .I1(\trig_pc_reg[63]_0 [6]),
        .I2(\wb_reg_pc_reg[39]_0 [6]),
        .I3(\trig_pc_reg[63]_0 [7]),
        .I4(\trig_pc_reg[63]_0 [8]),
        .I5(\wb_reg_pc_reg[39]_0 [7]),
        .O(\trig_pc_reg[0]_2 [2]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    core__266_i_28
       (.I0(\wb_reg_pc_reg[39]_0 [2]),
        .I1(\trig_pc_reg[63]_0 [3]),
        .I2(\wb_reg_pc_reg[39]_0 [3]),
        .I3(\trig_pc_reg[63]_0 [4]),
        .I4(\trig_pc_reg[63]_0 [5]),
        .I5(\wb_reg_pc_reg[39]_0 [4]),
        .O(\trig_pc_reg[0]_2 [1]));
  LUT5 #(
    .INIT(32'h41000041)) 
    core__266_i_29
       (.I0(\trig_pc_reg[63]_0 [0]),
        .I1(\wb_reg_pc_reg[39]_0 [0]),
        .I2(\trig_pc_reg[63]_0 [1]),
        .I3(\trig_pc_reg[63]_0 [2]),
        .I4(\wb_reg_pc_reg[39]_0 [1]),
        .O(\trig_pc_reg[0]_2 [0]));
  LUT3 #(
    .INIT(8'h01)) 
    core__266_i_5
       (.I0(\trig_pc_reg[63]_0 [61]),
        .I1(\trig_pc_reg[63]_0 [60]),
        .I2(\trig_pc_reg[63]_0 [62]),
        .O(\trig_pc_reg[0]_7 ));
  LUT3 #(
    .INIT(8'h01)) 
    core__266_i_7
       (.I0(\trig_pc_reg[63]_0 [58]),
        .I1(\trig_pc_reg[63]_0 [57]),
        .I2(\trig_pc_reg[63]_0 [59]),
        .O(\trig_pc_reg[0]_6 [3]));
  LUT3 #(
    .INIT(8'h01)) 
    core__266_i_8
       (.I0(\trig_pc_reg[63]_0 [55]),
        .I1(\trig_pc_reg[63]_0 [54]),
        .I2(\trig_pc_reg[63]_0 [56]),
        .O(\trig_pc_reg[0]_6 [2]));
  LUT3 #(
    .INIT(8'h01)) 
    core__266_i_9
       (.I0(\trig_pc_reg[63]_0 [52]),
        .I1(\trig_pc_reg[63]_0 [51]),
        .I2(\trig_pc_reg[63]_0 [53]),
        .O(\trig_pc_reg[0]_6 [1]));
  (* SOFT_HLUTNM = "soft_lutpair1786" *) 
  LUT2 #(
    .INIT(4'hB)) 
    core__268_i_1
       (.I0(ex_ctrl_sel_alu2[0]),
        .I1(ex_ctrl_sel_alu2[1]),
        .O(\bypass_mux_1_reg[4]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1790" *) 
  LUT5 #(
    .INIT(32'h24FFFFFF)) 
    core__268_i_2
       (.I0(\bypass_mux_1_reg[6]_1 [2]),
        .I1(\bypass_mux_1_reg[6]_1 [1]),
        .I2(\bypass_mux_1_reg[6]_1 [0]),
        .I3(ex_ctrl_sel_alu2[1]),
        .I4(ex_ctrl_sel_alu2[0]),
        .O(\bypass_mux_1_reg[6]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1857" *) 
  LUT4 #(
    .INIT(16'h3404)) 
    core__292_i_1
       (.I0(neg_out_reg),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[39]),
        .O(alu_io_in1[62]));
  LUT4 #(
    .INIT(16'hFF40)) 
    core__292_i_2
       (.I0(ex_ctrl_sel_alu2[0]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(mem_reg_rs2[63]),
        .I3(\ex_ctrl_sel_imm_reg[1]_0 ),
        .O(alu_io_in2[62]));
  (* SOFT_HLUTNM = "soft_lutpair1789" *) 
  LUT4 #(
    .INIT(16'h0200)) 
    core__434_i_1
       (.I0(mem_ctrl_branch),
        .I1(\trig_state_reg[1]_0 ),
        .I2(\trig_state_reg[0]_0 ),
        .I3(\trig_state_reg[1]_1 ),
        .O(trig_pc_valid_reg_0));
  (* SOFT_HLUTNM = "soft_lutpair1826" *) 
  LUT3 #(
    .INIT(8'h08)) 
    core__434_i_2
       (.I0(\trig_state_reg[0]_0 ),
        .I1(\trig_state_reg[1]_0 ),
        .I2(\trig_state_reg[1]_1 ),
        .O(\trig_jalr_count_reg[0]_0 ));
  LUT4 #(
    .INIT(16'h3808)) 
    core__436_i_1
       (.I0(div_n_139),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[2]),
        .O(alu_io_in1[1]));
  LUT6 #(
    .INIT(64'h30FF550030005500)) 
    core__436_i_2
       (.I0(mem_reg_rvc_reg_0),
        .I1(core__168_i_5_n_0),
        .I2(core__436_i_3_n_0),
        .I3(ex_ctrl_sel_alu2[0]),
        .I4(ex_ctrl_sel_alu2[1]),
        .I5(mem_reg_rs2[2]),
        .O(alu_io_in2[2]));
  LUT6 #(
    .INIT(64'hFECEFEFE32020202)) 
    core__436_i_3
       (.I0(\mem_reg_inst_reg[31]_0 [2]),
        .I1(\bypass_mux_1_reg[6]_1 [1]),
        .I2(\bypass_mux_1_reg[6]_1 [2]),
        .I3(\ex_reg_inst_reg_n_0_[17] ),
        .I4(\bypass_mux_1_reg[6]_1 [0]),
        .I5(\ex_reg_inst_reg_n_0_[22] ),
        .O(core__436_i_3_n_0));
  LUT4 #(
    .INIT(16'h3808)) 
    core__439_i_1
       (.I0(div_n_142),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[5]),
        .O(alu_io_in1[4]));
  LUT5 #(
    .INIT(32'h40FF4040)) 
    core__439_i_2
       (.I0(ex_ctrl_sel_alu2[0]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(mem_reg_rs2[5]),
        .I3(\bypass_mux_1_reg[6]_0 ),
        .I4(\ex_reg_inst_reg_n_0_[25] ),
        .O(alu_io_in2[5]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__440_i_1
       (.I0(div_n_143),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[6]),
        .O(alu_io_in1[5]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__441_i_1
       (.I0(div_n_148),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[11]),
        .O(alu_io_in1[10]));
  (* SOFT_HLUTNM = "soft_lutpair1786" *) 
  LUT5 #(
    .INIT(32'h04FF0404)) 
    core__441_i_2
       (.I0(ex_ctrl_sel_alu2[0]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(div_n_220),
        .I3(\bypass_mux_1_reg[6]_0 ),
        .I4(core__441_i_3_n_0),
        .O(alu_io_in2[10]));
  LUT6 #(
    .INIT(64'hE3FFE0FF23002000)) 
    core__441_i_3
       (.I0(_T_1710),
        .I1(\bypass_mux_1_reg[6]_1 [2]),
        .I2(\bypass_mux_1_reg[6]_1 [1]),
        .I3(\bypass_mux_1_reg[6]_1 [0]),
        .I4(\mem_reg_inst_reg[31]_0 [0]),
        .I5(\mem_reg_inst_reg[31]_0 [7]),
        .O(core__441_i_3_n_0));
  LUT4 #(
    .INIT(16'h3808)) 
    core__442_i_1
       (.I0(div_n_149),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[12]),
        .O(alu_io_in1[11]));
  LUT6 #(
    .INIT(64'hC404C4C4C4040404)) 
    core__442_i_2
       (.I0(div_n_221),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[12] ),
        .I4(core__166_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[11]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__443_i_1
       (.I0(div_n_152),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[15]),
        .O(alu_io_in1[14]));
  LUT6 #(
    .INIT(64'hC404C4C4C4040404)) 
    core__443_i_2
       (.I0(div_n_224),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[15] ),
        .I4(core__166_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[14]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__444_i_1
       (.I0(div_n_155),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[18]),
        .O(alu_io_in1[17]));
  LUT6 #(
    .INIT(64'hC404C4C4C4040404)) 
    core__444_i_2
       (.I0(div_n_225),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[18] ),
        .I4(core__166_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[17]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__445_i_1
       (.I0(div_n_158),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[21]),
        .O(alu_io_in1[20]));
  LUT6 #(
    .INIT(64'hC404C4C4C4040404)) 
    core__445_i_2
       (.I0(div_n_228),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[21] ),
        .I4(core__168_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[20]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__446_i_1
       (.I0(div_n_161),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[24]),
        .O(alu_io_in1[23]));
  LUT6 #(
    .INIT(64'hC808C8C8C8080808)) 
    core__446_i_2
       (.I0(mem_reg_rs2[24]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[24] ),
        .I4(core__168_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[23]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__447_i_1
       (.I0(div_n_164),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[27]),
        .O(alu_io_in1[26]));
  LUT6 #(
    .INIT(64'hC808C8C8C8080808)) 
    core__447_i_2
       (.I0(mem_reg_rs2[27]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\mem_reg_inst_reg[31]_0 [6]),
        .I4(core__168_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[26]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__448_i_1
       (.I0(div_n_167),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[30]),
        .O(alu_io_in1[29]));
  LUT6 #(
    .INIT(64'hC808C8C8C8080808)) 
    core__448_i_2
       (.I0(mem_reg_rs2[30]),
        .I1(ex_ctrl_sel_alu2[1]),
        .I2(ex_ctrl_sel_alu2[0]),
        .I3(\ex_reg_inst_reg_n_0_[30] ),
        .I4(core__168_i_5_n_0),
        .I5(core__166_i_6_n_0),
        .O(alu_io_in2[29]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__449_i_1
       (.I0(\remainder_reg[33]_0 ),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[33]),
        .O(alu_io_in1[32]));
  (* SOFT_HLUTNM = "soft_lutpair1843" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__449_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[33]),
        .O(alu_io_in2[32]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__450_i_1
       (.I0(\remainder_reg[36]_0 ),
        .I1(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I3(ex_reg_pc[36]),
        .O(alu_io_in1[35]));
  (* SOFT_HLUTNM = "soft_lutpair1847" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__450_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[36]),
        .O(alu_io_in2[35]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__451_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [0]),
        .O(alu_io_in1[38]));
  (* SOFT_HLUTNM = "soft_lutpair1852" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__451_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[39]),
        .O(alu_io_in2[38]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__452_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [2]),
        .O(alu_io_in1[41]));
  (* SOFT_HLUTNM = "soft_lutpair1858" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__452_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[42]),
        .O(alu_io_in2[41]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__453_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(_T_2770[6]),
        .O(alu_io_in1[44]));
  (* SOFT_HLUTNM = "soft_lutpair1854" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__453_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[45]),
        .O(alu_io_in2[44]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__454_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(_T_2770[9]),
        .O(alu_io_in1[47]));
  (* SOFT_HLUTNM = "soft_lutpair1850" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__454_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[48]),
        .O(alu_io_in2[47]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__455_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [9]),
        .O(alu_io_in1[50]));
  (* SOFT_HLUTNM = "soft_lutpair1855" *) 
  LUT4 #(
    .INIT(16'hAABA)) 
    core__455_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(div_n_235),
        .O(alu_io_in2[50]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__456_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [11]),
        .O(alu_io_in1[53]));
  (* SOFT_HLUTNM = "soft_lutpair1861" *) 
  LUT4 #(
    .INIT(16'hAABA)) 
    core__456_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(div_n_238),
        .O(alu_io_in2[53]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__457_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [13]),
        .O(alu_io_in1[56]));
  (* SOFT_HLUTNM = "soft_lutpair1859" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__457_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(\divisor_reg[57] [5]),
        .O(alu_io_in2[56]));
  LUT4 #(
    .INIT(16'h3808)) 
    core__458_i_1
       (.I0(ex_reg_pc[39]),
        .I1(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .I2(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .I3(\s1_req_addr_reg[39] [15]),
        .O(alu_io_in1[59]));
  (* SOFT_HLUTNM = "soft_lutpair1843" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    core__458_i_2
       (.I0(\ex_ctrl_sel_imm_reg[1]_0 ),
        .I1(ex_ctrl_sel_alu2[0]),
        .I2(ex_ctrl_sel_alu2[1]),
        .I3(mem_reg_rs2[60]),
        .O(alu_io_in2[59]));
  LUT2 #(
    .INIT(4'h7)) 
    core__462_i_13
       (.I0(wb_reg_cause[63]),
        .I1(wb_reg_xcpt),
        .O(\reg_sbadaddr_reg[30]_9 [1]));
  LUT1 #(
    .INIT(2'h1)) 
    core__462_i_14
       (.I0(core__506_i_2_n_0),
        .O(\reg_sbadaddr_reg[30]_9 [0]));
  LUT2 #(
    .INIT(4'h7)) 
    core__462_i_15
       (.I0(wb_reg_cause[63]),
        .I1(wb_reg_xcpt),
        .O(\reg_sbadaddr_reg[30]_1 [2]));
  LUT1 #(
    .INIT(2'h1)) 
    core__462_i_16
       (.I0(core__506_i_2_n_0),
        .O(\reg_sbadaddr_reg[30]_1 [1]));
  LUT4 #(
    .INIT(16'h0004)) 
    core__462_i_17
       (.I0(\reg_scause_reg[1] ),
        .I1(wb_reg_xcpt),
        .I2(\reg_scause_reg[2] ),
        .I3(\reg_scause_reg[0]_0 ),
        .O(\reg_sbadaddr_reg[30]_1 [0]));
  LUT2 #(
    .INIT(4'h7)) 
    core__462_i_18
       (.I0(wb_reg_cause[63]),
        .I1(wb_reg_xcpt),
        .O(\reg_sbadaddr_reg[30]_6 [2]));
  LUT6 #(
    .INIT(64'hFF000000FF0EFF0E)) 
    core__462_i_19
       (.I0(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
        .I1(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
        .I2(\lrscCount_reg[0] ),
        .I3(wb_reg_xcpt),
        .I4(wb_reg_cause[3]),
        .I5(\lrscCount_reg[0]_0 ),
        .O(\reg_sbadaddr_reg[30]_6 [1]));
  LUT4 #(
    .INIT(16'h00A2)) 
    core__462_i_20
       (.I0(\reg_scause_reg[0]_0 ),
        .I1(wb_reg_xcpt),
        .I2(\reg_scause_reg[2] ),
        .I3(\reg_scause_reg[1] ),
        .O(\reg_sbadaddr_reg[30]_6 [0]));
  LUT2 #(
    .INIT(4'h7)) 
    core__462_i_21
       (.I0(wb_reg_cause[63]),
        .I1(wb_reg_xcpt),
        .O(\reg_sbadaddr_reg[30] [2]));
  LUT1 #(
    .INIT(2'h1)) 
    core__462_i_22
       (.I0(core__506_i_2_n_0),
        .O(\reg_sbadaddr_reg[30] [1]));
  LUT4 #(
    .INIT(16'h8808)) 
    core__462_i_23
       (.I0(\reg_scause_reg[0]_0 ),
        .I1(\reg_scause_reg[1] ),
        .I2(wb_reg_xcpt),
        .I3(\reg_scause_reg[2] ),
        .O(\reg_sbadaddr_reg[30] [0]));
  LUT2 #(
    .INIT(4'h7)) 
    core__462_i_24
       (.I0(wb_reg_cause[63]),
        .I1(wb_reg_xcpt),
        .O(\reg_sbadaddr_reg[30]_0 [2]));
  LUT1 #(
    .INIT(2'h1)) 
    core__462_i_25
       (.I0(core__506_i_2_n_0),
        .O(\reg_sbadaddr_reg[30]_0 [1]));
  LUT4 #(
    .INIT(16'h0008)) 
    core__462_i_26
       (.I0(\reg_scause_reg[1] ),
        .I1(wb_reg_xcpt),
        .I2(\reg_scause_reg[2] ),
        .I3(\reg_scause_reg[0]_0 ),
        .O(\reg_sbadaddr_reg[30]_0 [0]));
  LUT2 #(
    .INIT(4'h7)) 
    core__462_i_27
       (.I0(wb_reg_cause[63]),
        .I1(wb_reg_xcpt),
        .O(\reg_sbadaddr_reg[30]_2 [1]));
  LUT1 #(
    .INIT(2'h1)) 
    core__462_i_28
       (.I0(core__506_i_2_n_0),
        .O(\reg_sbadaddr_reg[30]_2 [0]));
  LUT2 #(
    .INIT(4'h7)) 
    core__462_i_29
       (.I0(wb_reg_cause[63]),
        .I1(wb_reg_xcpt),
        .O(\reg_sbadaddr_reg[30]_4 [2]));
  LUT1 #(
    .INIT(2'h1)) 
    core__462_i_30
       (.I0(core__506_i_2_n_0),
        .O(\reg_sbadaddr_reg[30]_4 [1]));
  LUT4 #(
    .INIT(16'h00A2)) 
    core__462_i_31
       (.I0(\reg_scause_reg[0]_0 ),
        .I1(wb_reg_xcpt),
        .I2(\reg_scause_reg[2] ),
        .I3(\reg_scause_reg[1] ),
        .O(\reg_sbadaddr_reg[30]_4 [0]));
  LUT2 #(
    .INIT(4'h7)) 
    core__462_i_32
       (.I0(wb_reg_cause[63]),
        .I1(wb_reg_xcpt),
        .O(\reg_sbadaddr_reg[30]_8 [1]));
  LUT6 #(
    .INIT(64'hFF000000FF0EFF0E)) 
    core__462_i_33
       (.I0(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
        .I1(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
        .I2(\lrscCount_reg[0] ),
        .I3(wb_reg_xcpt),
        .I4(wb_reg_cause[3]),
        .I5(\lrscCount_reg[0]_0 ),
        .O(\reg_sbadaddr_reg[30]_8 [0]));
  LUT2 #(
    .INIT(4'h7)) 
    core__462_i_34
       (.I0(wb_reg_cause[63]),
        .I1(wb_reg_xcpt),
        .O(\reg_sbadaddr_reg[30]_7 [1]));
  LUT6 #(
    .INIT(64'hFF000000FF0EFF0E)) 
    core__462_i_35
       (.I0(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
        .I1(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
        .I2(\lrscCount_reg[0] ),
        .I3(wb_reg_xcpt),
        .I4(wb_reg_cause[3]),
        .I5(\lrscCount_reg[0]_0 ),
        .O(\reg_sbadaddr_reg[30]_7 [0]));
  LUT2 #(
    .INIT(4'h7)) 
    core__462_i_36
       (.I0(wb_reg_cause[63]),
        .I1(wb_reg_xcpt),
        .O(\reg_sbadaddr_reg[30]_5 [1]));
  LUT1 #(
    .INIT(2'h1)) 
    core__462_i_37
       (.I0(core__506_i_2_n_0),
        .O(\reg_sbadaddr_reg[30]_5 [0]));
  (* SOFT_HLUTNM = "soft_lutpair1867" *) 
  LUT3 #(
    .INIT(8'h08)) 
    core__49_i_1
       (.I0(ex_ctrl_wxd),
        .I1(ex_reg_valid),
        .I2(\ex_reg_inst_reg[10]_0 ),
        .O(\ex_reg_rs_lsb_0_reg[0]_1 ));
  LUT3 #(
    .INIT(8'hFD)) 
    core__4_i_1
       (.I0(\ex_reg_rs_lsb_0_reg[0]_0 ),
        .I1(\ex_reg_rs_lsb_0_reg[0]_1 ),
        .I2(nBufValid_reg_5),
        .O(_T_1829));
  (* SOFT_HLUTNM = "soft_lutpair1821" *) 
  LUT5 #(
    .INIT(32'h0010FFFE)) 
    core__506_i_1
       (.I0(\wb_ctrl_csr_reg[0]_0 ),
        .I1(\reg_bp_0_control_tmatch_reg[1] [6]),
        .I2(\reg_bp_0_control_tmatch_reg[1] [5]),
        .I3(\reg_bp_0_control_tmatch_reg[1] [7]),
        .I4(core__506_i_2_n_0),
        .O(\reg_scause_reg[3] ));
  LUT6 #(
    .INIT(64'hFF000000FF0EFF0E)) 
    core__506_i_2
       (.I0(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
        .I1(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
        .I2(\lrscCount_reg[0] ),
        .I3(wb_reg_xcpt),
        .I4(wb_reg_cause[3]),
        .I5(\lrscCount_reg[0]_0 ),
        .O(core__506_i_2_n_0));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__638_i_1
       (.I0(\bypass_mux_1_reg[33]_3 ),
        .I1(\bypass_mux_1_reg[38]_2 ),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[33]_4 ),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[42]_2 ),
        .O(\bypass_mux_1_reg[33]_2 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__638_i_2
       (.I0(core__638_i_4_n_0),
        .I1(\bypass_mux_1_reg[40]_2 ),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[35]_3 ),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[44]_2 ),
        .O(\bypass_mux_1_reg[35]_2 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__638_i_3
       (.I0(\bypass_mux_1_reg[34]_3 ),
        .I1(\bypass_mux_1_reg[39]_2 ),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[34]_4 ),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[43]_2 ),
        .O(\bypass_mux_1_reg[34]_2 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__638_i_4
       (.I0(\alu/shin [59]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [43]),
        .O(core__638_i_4_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1792" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__638_i_5
       (.I0(alu_io_in1[58]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[3]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [59]));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__639_i_1
       (.I0(\alu/shin [55]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [39]),
        .O(\bypass_mux_1_reg[35]_3 ));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__639_i_10
       (.I0(\alu/shin [59]),
        .I1(shamt),
        .I2(alu_io_in1[26]),
        .I3(core__639_i_11_n_0),
        .I4(\alu/_T_55 ),
        .O(core__639_i_10_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1813" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__639_i_11
       (.I0(alu_io_in1[35]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__639_i_11_n_0));
  LUT6 #(
    .INIT(64'hAF00CFCFAF00C0C0)) 
    core__639_i_2
       (.I0(Q),
        .I1(\bypass_mux_1_reg[1]_0 [2]),
        .I2(alu_io_in2[4]),
        .I3(\bypass_mux_1_reg[1]_0 [3]),
        .I4(shamt),
        .I5(\bypass_mux_1_reg[1]_0 [1]),
        .O(\bypass_mux_1_reg[44]_2 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__639_i_3
       (.I0(\alu/shin [51]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [35]),
        .O(\bypass_mux_1_reg[40]_2 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__639_i_4
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [43]),
        .I3(alu_io_in2[4]),
        .I4(core__639_i_10_n_0),
        .O(\bypass_mux_1_reg[48]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair1796" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__639_i_5
       (.I0(alu_io_in1[54]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[7]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [55]));
  (* SOFT_HLUTNM = "soft_lutpair1809" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__639_i_6
       (.I0(alu_io_in1[38]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[23]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [39]));
  (* SOFT_HLUTNM = "soft_lutpair1800" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__639_i_7
       (.I0(alu_io_in1[50]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[11]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [51]));
  (* SOFT_HLUTNM = "soft_lutpair1817" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__639_i_8
       (.I0(alu_io_in1[34]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[27]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [35]));
  (* SOFT_HLUTNM = "soft_lutpair1805" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__639_i_9
       (.I0(alu_io_in1[42]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[19]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [43]));
  (* SOFT_HLUTNM = "soft_lutpair1840" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__640_i_1
       (.I0(alu_io_in1[62]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(\bypass_mux_1_reg[0]_0 ),
        .I4(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[1]_0 [3]));
  LUT2 #(
    .INIT(4'h8)) 
    core__640_i_2
       (.I0(alu_io_in2[5]),
        .I1(req_dw_reg),
        .O(shamt));
  (* SOFT_HLUTNM = "soft_lutpair1819" *) 
  LUT5 #(
    .INIT(32'hF0F0B888)) 
    core__640_i_3
       (.I0(alu_io_in1[31]),
        .I1(req_dw_reg),
        .I2(alu_io_in1[30]),
        .I3(Q),
        .I4(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[1]_0 [1]));
  (* SOFT_HLUTNM = "soft_lutpair1804" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__640_i_4
       (.I0(alu_io_in1[46]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[15]),
        .I4(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[1]_0 [2]));
  (* SOFT_HLUTNM = "soft_lutpair1803" *) 
  LUT5 #(
    .INIT(32'hAAAACFC0)) 
    core__640_i_5
       (.I0(alu_io_in1[14]),
        .I1(alu_io_in1[47]),
        .I2(req_dw_reg),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(\alu/_T_55 ),
        .O(\bypass_mux_1_reg[1]_0 [0]));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__641_i_1
       (.I0(\alu/shin [56]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [40]),
        .O(\bypass_mux_1_reg[34]_4 ));
  (* SOFT_HLUTNM = "soft_lutpair1813" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__641_i_10
       (.I0(alu_io_in1[35]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[26]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [36]));
  (* SOFT_HLUTNM = "soft_lutpair1808" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__641_i_11
       (.I0(alu_io_in1[43]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[18]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [44]));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__641_i_12
       (.I0(\alu/shin [60]),
        .I1(shamt),
        .I2(alu_io_in1[27]),
        .I3(core__641_i_13_n_0),
        .I4(\alu/_T_55 ),
        .O(core__641_i_12_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1817" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__641_i_13
       (.I0(alu_io_in1[34]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__641_i_13_n_0));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__641_i_2
       (.I0(\alu/shin [48]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [32]),
        .O(\bypass_mux_1_reg[43]_2 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__641_i_3
       (.I0(\alu/shin [52]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [36]),
        .O(\bypass_mux_1_reg[39]_2 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__641_i_4
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [44]),
        .I3(alu_io_in2[4]),
        .I4(core__641_i_12_n_0),
        .O(\bypass_mux_1_reg[47]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair1795" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__641_i_5
       (.I0(alu_io_in1[55]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[6]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [56]));
  (* SOFT_HLUTNM = "soft_lutpair1812" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__641_i_6
       (.I0(alu_io_in1[39]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[22]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [40]));
  (* SOFT_HLUTNM = "soft_lutpair1803" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__641_i_7
       (.I0(alu_io_in1[47]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[14]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [48]));
  (* SOFT_HLUTNM = "soft_lutpair1819" *) 
  LUT5 #(
    .INIT(32'hF8AA08AA)) 
    core__641_i_8
       (.I0(alu_io_in1[30]),
        .I1(Q),
        .I2(req_dw_reg),
        .I3(\alu/_T_55 ),
        .I4(alu_io_in1[31]),
        .O(\alu/shin [32]));
  (* SOFT_HLUTNM = "soft_lutpair1799" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__641_i_9
       (.I0(alu_io_in1[51]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[10]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [52]));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__642_i_1
       (.I0(\bypass_mux_1_reg[29]_4 ),
        .I1(\bypass_mux_1_reg[35]_3 ),
        .I2(alu_io_in2[2]),
        .I3(core__638_i_4_n_0),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[40]_2 ),
        .O(\bypass_mux_1_reg[29]_1 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    core__642_i_2
       (.I0(\bypass_mux_1_reg[29]_2 ),
        .I1(\bypass_mux_1_reg[37]_2 ),
        .I2(alu_io_in2[2]),
        .I3(\bypass_mux_1_reg[29]_3 ),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[41]_2 ),
        .O(\bypass_mux_1_reg[29]_0 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__643_i_1
       (.I0(\alu/shin [57]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [41]),
        .O(\bypass_mux_1_reg[33]_4 ));
  (* SOFT_HLUTNM = "soft_lutpair1816" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__643_i_10
       (.I0(alu_io_in1[36]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[25]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [37]));
  (* SOFT_HLUTNM = "soft_lutpair1807" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__643_i_11
       (.I0(alu_io_in1[44]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[17]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [45]));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__643_i_12
       (.I0(\alu/shin [61]),
        .I1(shamt),
        .I2(alu_io_in1[28]),
        .I3(core__643_i_13_n_0),
        .I4(\alu/_T_55 ),
        .O(core__643_i_12_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1818" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__643_i_13
       (.I0(alu_io_in1[33]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__643_i_13_n_0));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__643_i_2
       (.I0(\alu/shin [49]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [33]),
        .O(\bypass_mux_1_reg[42]_2 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__643_i_3
       (.I0(\alu/shin [53]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [37]),
        .O(\bypass_mux_1_reg[38]_2 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__643_i_4
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [45]),
        .I3(alu_io_in2[4]),
        .I4(core__643_i_12_n_0),
        .O(\bypass_mux_1_reg[46]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair1794" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__643_i_5
       (.I0(alu_io_in1[56]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[5]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [57]));
  (* SOFT_HLUTNM = "soft_lutpair1810" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__643_i_6
       (.I0(alu_io_in1[40]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[21]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [41]));
  (* SOFT_HLUTNM = "soft_lutpair1785" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__643_i_7
       (.I0(alu_io_in1[48]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[13]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [49]));
  (* SOFT_HLUTNM = "soft_lutpair1820" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__643_i_8
       (.I0(alu_io_in1[32]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[29]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [33]));
  (* SOFT_HLUTNM = "soft_lutpair1798" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__643_i_9
       (.I0(alu_io_in1[52]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[9]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [53]));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__644_i_1
       (.I0(\alu/shin [58]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [42]),
        .O(\bypass_mux_1_reg[29]_3 ));
  (* SOFT_HLUTNM = "soft_lutpair1815" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__644_i_10
       (.I0(alu_io_in1[37]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[24]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [38]));
  (* SOFT_HLUTNM = "soft_lutpair1806" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__644_i_11
       (.I0(alu_io_in1[45]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[16]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [46]));
  LUT5 #(
    .INIT(32'hB8B8BB88)) 
    core__644_i_12
       (.I0(\alu/shin [62]),
        .I1(shamt),
        .I2(alu_io_in1[29]),
        .I3(core__644_i_13_n_0),
        .I4(\alu/_T_55 ),
        .O(core__644_i_12_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1820" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__644_i_13
       (.I0(alu_io_in1[32]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .O(core__644_i_13_n_0));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__644_i_2
       (.I0(\alu/shin [50]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [34]),
        .O(\bypass_mux_1_reg[41]_2 ));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__644_i_3
       (.I0(\alu/shin [54]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [38]),
        .O(\bypass_mux_1_reg[37]_2 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    core__644_i_4
       (.I0(_T_121),
        .I1(shamt),
        .I2(\alu/shin [46]),
        .I3(alu_io_in2[4]),
        .I4(core__644_i_12_n_0),
        .O(\bypass_mux_1_reg[45]_2 ));
  (* SOFT_HLUTNM = "soft_lutpair1793" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__644_i_5
       (.I0(alu_io_in1[57]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[4]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [58]));
  (* SOFT_HLUTNM = "soft_lutpair1811" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__644_i_6
       (.I0(alu_io_in1[41]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[20]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [42]));
  (* SOFT_HLUTNM = "soft_lutpair1801" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__644_i_7
       (.I0(alu_io_in1[49]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[12]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [50]));
  (* SOFT_HLUTNM = "soft_lutpair1818" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__644_i_8
       (.I0(alu_io_in1[33]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[28]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [34]));
  (* SOFT_HLUTNM = "soft_lutpair1797" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__644_i_9
       (.I0(alu_io_in1[53]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[8]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [54]));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__645_i_1
       (.I0(\alu/shin [60]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [44]),
        .O(\bypass_mux_1_reg[34]_3 ));
  LUT6 #(
    .INIT(64'hCDC8FFFFCDC80000)) 
    core__645_i_2
       (.I0(alu_io_in2[4]),
        .I1(_T_121),
        .I2(shamt),
        .I3(\alu/shin [48]),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[34]_4 ),
        .O(\bypass_mux_1_reg[23]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1788" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__645_i_3
       (.I0(alu_io_in1[59]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[2]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [60]));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__646_i_1
       (.I0(\alu/shin [61]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [45]),
        .O(\bypass_mux_1_reg[33]_3 ));
  LUT6 #(
    .INIT(64'hCDC8FFFFCDC80000)) 
    core__646_i_2
       (.I0(alu_io_in2[4]),
        .I1(_T_121),
        .I2(shamt),
        .I3(\alu/shin [49]),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[33]_4 ),
        .O(\bypass_mux_1_reg[22]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1784" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__646_i_3
       (.I0(alu_io_in1[60]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[1]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [61]));
  LUT5 #(
    .INIT(32'hF0BBF088)) 
    core__647_i_1
       (.I0(\alu/shin [62]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [46]),
        .O(\bypass_mux_1_reg[29]_2 ));
  LUT6 #(
    .INIT(64'hCDC8FFFFCDC80000)) 
    core__647_i_2
       (.I0(alu_io_in2[4]),
        .I1(_T_121),
        .I2(shamt),
        .I3(\alu/shin [50]),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[29]_3 ),
        .O(\bypass_mux_1_reg[21]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1791" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    core__647_i_3
       (.I0(alu_io_in1[61]),
        .I1(req_dw_reg),
        .I2(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I3(alu_io_in1[0]),
        .I4(\alu/_T_55 ),
        .O(\alu/shin [62]));
  LUT5 #(
    .INIT(32'hC0F5C0A0)) 
    core__648_i_1
       (.I0(alu_io_in2[4]),
        .I1(Q),
        .I2(\bypass_mux_1_reg[1]_0 [3]),
        .I3(shamt),
        .I4(\bypass_mux_1_reg[1]_0 [2]),
        .O(\bypass_mux_1_reg[29]_4 ));
  LUT6 #(
    .INIT(64'hCDC8FFFFCDC80000)) 
    core__648_i_2
       (.I0(alu_io_in2[4]),
        .I1(_T_121),
        .I2(shamt),
        .I3(\alu/shin [51]),
        .I4(alu_io_in2[3]),
        .I5(core__638_i_4_n_0),
        .O(\bypass_mux_1_reg[20]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1870" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__649_i_1
       (.I0(core__649_i_5_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__649_i_6_n_0),
        .O(\bypass_mux_1_reg[50]_2 ));
  LUT6 #(
    .INIT(64'hFF00FB0BFF00F808)) 
    core__649_i_10
       (.I0(\alu/shin [57]),
        .I1(alu_io_in2[3]),
        .I2(alu_io_in2[4]),
        .I3(_T_121),
        .I4(shamt),
        .I5(\alu/shin [49]),
        .O(core__649_i_10_n_0));
  LUT6 #(
    .INIT(64'hFF00FB0BFF00F808)) 
    core__649_i_11
       (.I0(\alu/shin [59]),
        .I1(alu_io_in2[3]),
        .I2(alu_io_in2[4]),
        .I3(_T_121),
        .I4(shamt),
        .I5(\alu/shin [51]),
        .O(core__649_i_11_n_0));
  LUT6 #(
    .INIT(64'hCDC8FFFFCDC80000)) 
    core__649_i_12
       (.I0(alu_io_in2[4]),
        .I1(_T_121),
        .I2(shamt),
        .I3(\alu/shin [55]),
        .I4(alu_io_in2[3]),
        .I5(\bypass_mux_1_reg[29]_4 ),
        .O(core__649_i_12_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1865" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__649_i_2
       (.I0(core__649_i_7_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__649_i_8_n_0),
        .O(\bypass_mux_1_reg[18]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1869" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__649_i_3
       (.I0(core__649_i_9_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__649_i_10_n_0),
        .O(\bypass_mux_1_reg[17]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1873" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__649_i_4
       (.I0(core__649_i_11_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__649_i_12_n_0),
        .O(\bypass_mux_1_reg[19]_0 ));
  LUT6 #(
    .INIT(64'hFF00FB0BFF00F808)) 
    core__649_i_5
       (.I0(\alu/shin [62]),
        .I1(alu_io_in2[3]),
        .I2(alu_io_in2[4]),
        .I3(_T_121),
        .I4(shamt),
        .I5(\alu/shin [54]),
        .O(core__649_i_5_n_0));
  LUT6 #(
    .INIT(64'hFF00FB0BFF00F808)) 
    core__649_i_6
       (.I0(\alu/shin [58]),
        .I1(alu_io_in2[3]),
        .I2(alu_io_in2[4]),
        .I3(_T_121),
        .I4(shamt),
        .I5(\alu/shin [50]),
        .O(core__649_i_6_n_0));
  LUT6 #(
    .INIT(64'hFF00FB0BFF00F808)) 
    core__649_i_7
       (.I0(\alu/shin [60]),
        .I1(alu_io_in2[3]),
        .I2(alu_io_in2[4]),
        .I3(_T_121),
        .I4(shamt),
        .I5(\alu/shin [52]),
        .O(core__649_i_7_n_0));
  LUT6 #(
    .INIT(64'hFF00FB0BFF00F808)) 
    core__649_i_8
       (.I0(\alu/shin [56]),
        .I1(alu_io_in2[3]),
        .I2(alu_io_in2[4]),
        .I3(_T_121),
        .I4(shamt),
        .I5(\alu/shin [48]),
        .O(core__649_i_8_n_0));
  LUT6 #(
    .INIT(64'hFF00FB0BFF00F808)) 
    core__649_i_9
       (.I0(\alu/shin [61]),
        .I1(alu_io_in2[3]),
        .I2(alu_io_in2[4]),
        .I3(_T_121),
        .I4(shamt),
        .I5(\alu/shin [53]),
        .O(core__649_i_9_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1871" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__650_i_1
       (.I0(core__650_i_2_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__649_i_11_n_0),
        .O(\bypass_mux_1_reg[51]_2 ));
  LUT6 #(
    .INIT(64'hF000F311F000E200)) 
    core__650_i_2
       (.I0(alu_io_in2[3]),
        .I1(alu_io_in2[4]),
        .I2(Q),
        .I3(\bypass_mux_1_reg[1]_0 [3]),
        .I4(shamt),
        .I5(\alu/shin [55]),
        .O(core__650_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1865" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__651_i_1
       (.I0(core__651_i_2_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__649_i_7_n_0),
        .O(\bypass_mux_1_reg[52]_2 ));
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    core__651_i_2
       (.I0(alu_io_in2[3]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [56]),
        .O(core__651_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1869" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__652_i_1
       (.I0(core__652_i_2_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__649_i_9_n_0),
        .O(\bypass_mux_1_reg[53]_2 ));
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    core__652_i_2
       (.I0(alu_io_in2[3]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [57]),
        .O(core__652_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1868" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__653_i_1
       (.I0(core__653_i_2_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__649_i_5_n_0),
        .O(\bypass_mux_1_reg[54]_2 ));
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    core__653_i_2
       (.I0(alu_io_in2[3]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [58]),
        .O(core__653_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1871" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__654_i_1
       (.I0(core__654_i_2_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__650_i_2_n_0),
        .O(\bypass_mux_1_reg[55]_2 ));
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    core__654_i_2
       (.I0(alu_io_in2[3]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [59]),
        .O(core__654_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1866" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__655_i_1
       (.I0(core__655_i_2_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__651_i_2_n_0),
        .O(\bypass_mux_1_reg[56]_2 ));
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    core__655_i_2
       (.I0(alu_io_in2[3]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [60]),
        .O(core__655_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1878" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__656_i_1
       (.I0(core__656_i_2_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__652_i_2_n_0),
        .O(\bypass_mux_1_reg[57]_2 ));
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    core__656_i_2
       (.I0(alu_io_in2[3]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [61]),
        .O(core__656_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1868" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__657_i_1
       (.I0(core__657_i_2_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__653_i_2_n_0),
        .O(\bypass_mux_1_reg[58]_2 ));
  LUT5 #(
    .INIT(32'hF0F1F0E0)) 
    core__657_i_2
       (.I0(alu_io_in2[3]),
        .I1(alu_io_in2[4]),
        .I2(_T_121),
        .I3(shamt),
        .I4(\alu/shin [62]),
        .O(core__657_i_2_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1875" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    core__658_i_1
       (.I0(core__658_i_2_n_0),
        .I1(alu_io_in2[2]),
        .I2(core__654_i_2_n_0),
        .O(\bypass_mux_1_reg[59]_2 ));
  LUT5 #(
    .INIT(32'hF0F10000)) 
    core__658_i_2
       (.I0(alu_io_in2[3]),
        .I1(alu_io_in2[4]),
        .I2(Q),
        .I3(shamt),
        .I4(\bypass_mux_1_reg[1]_0 [3]),
        .O(core__658_i_2_n_0));
  LUT6 #(
    .INIT(64'hFF00FF01FF00FE00)) 
    core__659_i_1
       (.I0(alu_io_in2[2]),
        .I1(alu_io_in2[3]),
        .I2(alu_io_in2[4]),
        .I3(_T_121),
        .I4(shamt),
        .I5(\alu/shin [60]),
        .O(\bypass_mux_1_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFF00FF01FF00FE00)) 
    core__660_i_1
       (.I0(alu_io_in2[2]),
        .I1(alu_io_in2[3]),
        .I2(alu_io_in2[4]),
        .I3(_T_121),
        .I4(shamt),
        .I5(\alu/shin [61]),
        .O(\bypass_mux_1_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFF00FF01FF00FE00)) 
    core__661_i_1
       (.I0(alu_io_in2[2]),
        .I1(alu_io_in2[3]),
        .I2(alu_io_in2[4]),
        .I3(_T_121),
        .I4(shamt),
        .I5(\alu/shin [62]),
        .O(\bypass_mux_1_reg[1]_2 ));
  LUT6 #(
    .INIT(64'hFF00FF0100000000)) 
    core__662_i_1
       (.I0(alu_io_in2[2]),
        .I1(alu_io_in2[3]),
        .I2(alu_io_in2[4]),
        .I3(Q),
        .I4(shamt),
        .I5(\bypass_mux_1_reg[1]_0 [3]),
        .O(\bypass_mux_1_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hA8A8A8202020A820)) 
    core__663_i_1
       (.I0(Q),
        .I1(\alu/_T_55 ),
        .I2(\bypass_mux_1_reg[0]_0 ),
        .I3(\ex_ctrl_alu_fn_reg[3]_8 ),
        .I4(req_dw_reg),
        .I5(alu_io_in1[62]),
        .O(_T_121));
  LUT6 #(
    .INIT(64'hFF2AFFFFFFFFFFFF)) 
    core__707_i_1
       (.I0(mem_reg_valid),
        .I1(core__707_i_3_n_0),
        .I2(core__707_i_4_n_0),
        .I3(wb_reg_flush_pipe),
        .I4(wb_reg_replay_reg_1),
        .I5(wb_reg_xcpt_i_2_n_0),
        .O(mem_reg_replay_reg_0));
  (* SOFT_HLUTNM = "soft_lutpair1862" *) 
  LUT2 #(
    .INIT(4'h1)) 
    core__707_i_3
       (.I0(mem_reg_sfence),
        .I1(mem_ctrl_jalr),
        .O(core__707_i_3_n_0));
  LUT6 #(
    .INIT(64'h1114111155555555)) 
    core__707_i_4
       (.I0(mem_ctrl_jal),
        .I1(mem_br_taken_),
        .I2(\trig_state_reg[1]_0 ),
        .I3(\trig_state_reg[0]_0 ),
        .I4(\trig_state_reg[1]_1 ),
        .I5(mem_ctrl_branch),
        .O(core__707_i_4_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    core__710_i_1
       (.I0(\trig_pc_reg[0]_0 ),
        .I1(\trig_pc_reg[63]_1 ),
        .O(\trig_state_reg[1]_2 ));
  CSRFile csr
       (.D({_T_5044[5],_T_5074,_T_4899,_T_5044[4:0]}),
        .Q(\reg_mtvec_reg[29] ),
        ._GEN_6(\bpu/_GEN_6 ),
        ._T_1005(_T_1005[0]),
        ._T_1081(_T_1081),
        ._T_1156(_T_1156),
        ._T_1432(_T_1432),
        ._T_1701(_T_1701),
        .\_T_1883_reg[0]_0 (\_T_1883_reg[0] ),
        .\_T_1883_reg[1]_0 (csr_io_status_debug),
        .\_T_1883_reg[1]_1 (\_T_1883_reg[1] ),
        ._T_200__0(_T_200__0),
        ._T_2177(_T_2177),
        ._T_2377(_T_2377),
        ._T_2518(_T_2518),
        .\_T_281_reg[0]_0 (\_T_281_reg[0] ),
        .\_T_281_reg[3]_0 (\_T_281_reg[3] ),
        .\_T_294_reg[0]_0 (\_T_294_reg[0] ),
        .\_T_294_reg[0]_1 (\_T_294_reg[0]_0 ),
        .\_T_294_reg[0]_2 (\_T_294_reg[0]_1 ),
        .\_T_294_reg[3]_0 (\_T_294_reg[3] ),
        ._T_382(_T_382),
        ._T_382_0(_T_382_0),
        ._T_382__0(_T_382__0),
        ._T_4068_ae_ld_reg(_T_4068_ae_ld_reg),
        ._T_4068_pf_ld_reg(_T_4068_pf_ld_reg),
        ._T_4068_pf_ld_reg_0(_T_4068_pf_ld_reg_0),
        ._T_4068_pf_ld_reg_1(_T_4068_pf_ld_reg_1),
        ._T_4068_pf_ld_reg_2(_T_4068_pf_ld_reg_2),
        ._T_4068_pf_ld_reg_3(_T_4068_pf_ld_reg_3),
        ._T_4068_pf_st_reg(_T_4068_pf_st_reg),
        ._T_4068_pf_st_reg_0(_T_4068_pf_st_reg_0),
        ._T_4068_pf_st_reg_1(_T_4068_pf_st_reg_1),
        ._T_480(_T_480),
        ._T_726(_T_726),
        ._T_931(_T_931),
        .\_T_973_reg[1] (\_T_973_reg[1] ),
        .bad_va(bad_va),
        .\buf__data_reg[12] (\buf__data_reg[12] ),
        .\buf__data_reg[3] (\buf__data_reg[3] ),
        .\buf__data_reg[3]_0 (\buf__data_reg[3]_0 ),
        .buf__xcpt_pf_inst_reg(buf__xcpt_pf_inst_reg),
        .buf__xcpt_pf_inst_reg_0(buf__xcpt_pf_inst_reg_0),
        .\bypass_mux_1_reg[32] ({\bypass_mux_1_reg_n_0_[32] ,\bypass_mux_1_reg_n_0_[31] ,\bypass_mux_1_reg_n_0_[30] ,\bypass_mux_1_reg_n_0_[29] ,\bypass_mux_1_reg_n_0_[28] ,\bypass_mux_1_reg_n_0_[27] ,\bypass_mux_1_reg_n_0_[26] ,\bypass_mux_1_reg_n_0_[25] ,\bypass_mux_1_reg_n_0_[24] ,\bypass_mux_1_reg_n_0_[23] ,\bypass_mux_1_reg_n_0_[22] ,\bypass_mux_1_reg_n_0_[21] ,\bypass_mux_1_reg_n_0_[20] ,\bypass_mux_1_reg_n_0_[19] ,\bypass_mux_1_reg_n_0_[18] ,\bypass_mux_1_reg_n_0_[17] ,\bypass_mux_1_reg_n_0_[16] ,\bypass_mux_1_reg_n_0_[15] ,\bypass_mux_1_reg_n_0_[14] ,\bypass_mux_1_reg_n_0_[13] ,\bypass_mux_1_reg_n_0_[12] ,\bypass_mux_1_reg_n_0_[11] ,\bypass_mux_1_reg_n_0_[10] ,\bypass_mux_1_reg_n_0_[9] ,\bypass_mux_1_reg_n_0_[8] ,\bypass_mux_1_reg_n_0_[7] ,\bypass_mux_1_reg_n_0_[6] ,\bypass_mux_1_reg_n_0_[5] ,\bypass_mux_1_reg_n_0_[4] ,\mem_reg_rs2_reg[3]_1 [1],\bypass_mux_1_reg_n_0_[2] ,\mem_reg_rs2_reg[3]_1 [0],\bypass_mux_1_reg_n_0_[0] }),
        .\bypass_mux_1_reg[33] (\bypass_mux_1_reg_n_0_[33] ),
        .\bypass_mux_1_reg[34] (\bypass_mux_1_reg_n_0_[34] ),
        .\bypass_mux_1_reg[35] (\bypass_mux_1_reg_n_0_[35] ),
        .\bypass_mux_1_reg[36] (\bypass_mux_1_reg_n_0_[36] ),
        .\bypass_mux_1_reg[36]_0 (\bypass_mux_1_reg[36]_2 ),
        .\bypass_mux_1_reg[37] (\bypass_mux_1_reg_n_0_[37] ),
        .\bypass_mux_1_reg[38] (\bypass_mux_2_reg[38]_0 ),
        .\bypass_mux_1_reg[38]_0 (\bypass_mux_1_reg[38]_3 ),
        .\bypass_mux_1_reg[39] (\s1_pc[39]_i_4_n_0 ),
        .\bypass_mux_2_reg[0] (\mem_reg_rs2_reg[0]_0 ),
        .\bypass_mux_2_reg[10] (\reg_mtvec_reg[10] ),
        .\bypass_mux_2_reg[11] (\reg_mtvec_reg[11] ),
        .\bypass_mux_2_reg[12] (\reg_mtvec_reg[12] ),
        .\bypass_mux_2_reg[13] (\reg_mtvec_reg[13] ),
        .\bypass_mux_2_reg[14] (\reg_mtvec_reg[14] ),
        .\bypass_mux_2_reg[15] (\reg_mtvec_reg[15] ),
        .\bypass_mux_2_reg[16] (\reg_mtvec_reg[16] ),
        .\bypass_mux_2_reg[17] (\reg_mtvec_reg[17] ),
        .\bypass_mux_2_reg[18] (\reg_mtvec_reg[18] ),
        .\bypass_mux_2_reg[19] (\reg_mtvec_reg[19] ),
        .\bypass_mux_2_reg[1] (\reg_misa_reg[12] [0]),
        .\bypass_mux_2_reg[1]_0 (\mem_reg_rs2_reg[1]_0 ),
        .\bypass_mux_2_reg[20] (\reg_mtvec_reg[20]_0 ),
        .\bypass_mux_2_reg[21] (\reg_mtvec_reg[21]_0 ),
        .\bypass_mux_2_reg[22] (\reg_mtvec_reg[22]_0 ),
        .\bypass_mux_2_reg[23] (\reg_mtvec_reg[23] ),
        .\bypass_mux_2_reg[24] (\reg_mtvec_reg[24] ),
        .\bypass_mux_2_reg[25] (\reg_mtvec_reg[25] ),
        .\bypass_mux_2_reg[26] (\reg_mtvec_reg[26] ),
        .\bypass_mux_2_reg[27] (\reg_mtvec_reg[27] ),
        .\bypass_mux_2_reg[28] (\reg_mtvec_reg[28] ),
        .\bypass_mux_2_reg[29] (\reg_mtvec_reg[29]_7 ),
        .\bypass_mux_2_reg[2] (\mem_reg_rs2_reg[2]_0 ),
        .\bypass_mux_2_reg[30] (\reg_mtvec_reg[30] ),
        .\bypass_mux_2_reg[31] (\reg_mtvec_reg[31] ),
        .\bypass_mux_2_reg[32] (\reg_stvec_reg[32] ),
        .\bypass_mux_2_reg[33] (\reg_stvec_reg[33] ),
        .\bypass_mux_2_reg[34] (\reg_stvec_reg[34] ),
        .\bypass_mux_2_reg[35] (\reg_stvec_reg[35] ),
        .\bypass_mux_2_reg[36] (\reg_stvec_reg[36] ),
        .\bypass_mux_2_reg[37] (\reg_stvec_reg[37] ),
        .\bypass_mux_2_reg[38] (\reg_stvec_reg[38] ),
        .\bypass_mux_2_reg[39] (\reg_sscratch_reg[62] [0]),
        .\bypass_mux_2_reg[3] (\mem_reg_rs2_reg[3]_0 ),
        .\bypass_mux_2_reg[40] (\reg_sscratch_reg[62] [1]),
        .\bypass_mux_2_reg[41] (\reg_sscratch_reg[62] [2]),
        .\bypass_mux_2_reg[42] (\reg_sscratch_reg[62] [3]),
        .\bypass_mux_2_reg[43] (\reg_sscratch_reg[62] [4]),
        .\bypass_mux_2_reg[44] (\reg_sscratch_reg[62] [5]),
        .\bypass_mux_2_reg[45] (\reg_sscratch_reg[62] [6]),
        .\bypass_mux_2_reg[46] (\reg_sscratch_reg[62] [7]),
        .\bypass_mux_2_reg[47] (\reg_sscratch_reg[62] [8]),
        .\bypass_mux_2_reg[48] (\reg_sscratch_reg[62] [9]),
        .\bypass_mux_2_reg[49] (\reg_sscratch_reg[62] [10]),
        .\bypass_mux_2_reg[4] (\mem_reg_rs2_reg[4]_0 ),
        .\bypass_mux_2_reg[50] (\reg_sscratch_reg[62] [11]),
        .\bypass_mux_2_reg[51] (\reg_sscratch_reg[62] [12]),
        .\bypass_mux_2_reg[52] (\reg_sscratch_reg[62] [13]),
        .\bypass_mux_2_reg[53] (\reg_sscratch_reg[62] [14]),
        .\bypass_mux_2_reg[54] (\reg_sscratch_reg[62] [15]),
        .\bypass_mux_2_reg[55] (\reg_sscratch_reg[62] [16]),
        .\bypass_mux_2_reg[56] (\reg_sscratch_reg[62] [17]),
        .\bypass_mux_2_reg[57] (\reg_sscratch_reg[62] [18]),
        .\bypass_mux_2_reg[58] (\reg_sscratch_reg[62] [19]),
        .\bypass_mux_2_reg[59] (\reg_sscratch_reg[62] [20]),
        .\bypass_mux_2_reg[5] (\mem_reg_rs2_reg[5]_0 ),
        .\bypass_mux_2_reg[60] (\reg_sscratch_reg[62] [21]),
        .\bypass_mux_2_reg[61] (\reg_sscratch_reg[62] [22]),
        .\bypass_mux_2_reg[62] (\reg_sscratch_reg[62] [23]),
        .\bypass_mux_2_reg[63] (\bypass_mux_2_reg[63]_0 ),
        .\bypass_mux_2_reg[63]_0 (\bypass_mux_2_reg[63]_1 ),
        .\bypass_mux_2_reg[6] (\mem_reg_rs2_reg[6]_0 ),
        .\bypass_mux_2_reg[7] (\mem_reg_rs2_reg[7]_0 ),
        .\bypass_mux_2_reg[8] (\reg_mtvec_reg[8] ),
        .\bypass_mux_2_reg[9] (reg_mip_seip_reg_0),
        .\count_reg[1] (\count_reg[1] ),
        .\count_reg[1]_0 (\count_reg[1]_0 ),
        .\count_reg[1]_1 (\count_reg[1]_1 ),
        .\count_reg[1]_2 (\count_reg[1]_2 ),
        .csr_io_bp_0_control_m(csr_io_bp_0_control_m),
        .csr_io_bp_0_control_s(csr_io_bp_0_control_s),
        .csr_io_bp_0_control_u(csr_io_bp_0_control_u),
        .csr_io_interrupt(csr_io_interrupt),
        .csr_io_tval(csr_io_tval),
        .dcacheArb_io_requestor_1_replay_next(dcacheArb_io_requestor_1_replay_next),
        .dcacheArb_io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),
        .dcacheArb_io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),
        .dcacheArb_io_requestor_1_s2_xcpt_ma_ld(dcacheArb_io_requestor_1_s2_xcpt_ma_ld),
        .dcacheArb_io_requestor_1_s2_xcpt_ma_st(dcacheArb_io_requestor_1_s2_xcpt_ma_st),
        .dcache_blocked(dcache_blocked),
        .dcache_io_cpu_invalidate_lr(dcache_io_cpu_invalidate_lr),
        .dcache_io_ptw_resp_bits_ae(dcache_io_ptw_resp_bits_ae),
        .dcache_io_ptw_resp_bits_homogeneous(dcache_io_ptw_resp_bits_homogeneous),
        .dcache_io_ptw_resp_bits_level(dcache_io_ptw_resp_bits_level),
        .dcache_io_ptw_resp_valid(dcache_io_ptw_resp_valid),
        .\elts_0_pc_reg[38] ({\elts_0_pc_reg[39] [17:16],ibuf_io_pc[36],\elts_0_pc_reg[39] [15],ibuf_io_pc[34],\elts_0_pc_reg[39] [14],ibuf_io_pc[32],\elts_0_pc_reg[39] [13],ibuf_io_pc[30],\elts_0_pc_reg[39] [12],ibuf_io_pc[28],\elts_0_pc_reg[39] [11],ibuf_io_pc[26],\elts_0_pc_reg[39] [10],ibuf_io_pc[24],\elts_0_pc_reg[39] [9],ibuf_io_pc[22],\elts_0_pc_reg[39] [8],ibuf_io_pc[20],\elts_0_pc_reg[39] [7],ibuf_io_pc[18],\elts_0_pc_reg[39] [6],ibuf_io_pc[16],\elts_0_pc_reg[39] [5],ibuf_io_pc[14],\elts_0_pc_reg[39] [4],ibuf_io_pc[12],\elts_0_pc_reg[39] [3],ibuf_io_pc[10],\elts_0_pc_reg[39] [2],ibuf_io_pc[8],\elts_0_pc_reg[39] [1],ibuf_io_pc[6],ibuf_io_pc[2:1]}),
        .\elts_0_pc_reg[38]_0 (\elts_0_pc_reg[38] ),
        .\ex_cause_reg[1] (\ex_cause_reg[1]_0 ),
        .\ex_cause_reg[1]_0 (_T_134),
        .\ex_cause_reg[1]_1 (\ex_cause_reg[1]_1 ),
        .\ex_cause_reg[1]_2 (\ex_cause_reg[1]_4 ),
        .\ex_cause_reg[1]_3 (\ex_cause_reg[1]_7 ),
        .\ex_cause_reg[1]_4 ({\ex_cause_reg[1]_12 [3:2],\ex_cause_reg[1]_12 [0]}),
        .\ex_cause_reg[3] ({csr_n_636,csr_n_637,csr_n_638,csr_n_639}),
        .\ex_cause_reg[63] (reg_dcsr_step),
        .\ex_cause_reg[63]_0 (reg_singleStepped),
        .ex_ctrl_div_reg(ex_ctrl_div),
        .ex_ctrl_mem_reg(ex_ctrl_mem_reg_0),
        .\ex_ctrl_sel_alu2_reg[1] (\ex_ctrl_sel_alu2_reg[1]_1 ),
        .\ex_ctrl_sel_alu2_reg[1]_0 (\ex_ctrl_sel_alu2_reg[1]_2 ),
        .\ex_ctrl_sel_alu2_reg[1]_1 (\ex_ctrl_sel_alu2_reg[1]_5 ),
        .\ex_ctrl_sel_alu2_reg[1]_2 (\ex_ctrl_sel_alu2_reg[1]_4 ),
        .\ex_reg_rs_lsb_1_reg[0] (csr_n_664),
        .\ex_reg_rs_lsb_1_reg[1] (csr_n_665),
        .\ex_reg_rs_msb_0_reg[10] (\ex_reg_rs_msb_0_reg[10]_0 ),
        .\ex_reg_rs_msb_0_reg[11] (\ex_reg_rs_msb_0_reg[11]_0 ),
        .\ex_reg_rs_msb_0_reg[12] (\ex_reg_rs_msb_0_reg[12]_0 ),
        .\ex_reg_rs_msb_0_reg[13] (\ex_reg_rs_msb_0_reg[13]_0 ),
        .\ex_reg_rs_msb_0_reg[14] (\ex_reg_rs_msb_0_reg[14]_0 ),
        .\ex_reg_rs_msb_0_reg[15] (\ex_reg_rs_msb_0_reg[15]_0 ),
        .\ex_reg_rs_msb_0_reg[16] (\ex_reg_rs_msb_0_reg[16]_0 ),
        .\ex_reg_rs_msb_0_reg[17] (\ex_reg_rs_msb_0_reg[17]_0 ),
        .\ex_reg_rs_msb_0_reg[18] (\ex_reg_rs_msb_0_reg[18]_0 ),
        .\ex_reg_rs_msb_0_reg[19] (\ex_reg_rs_msb_0_reg[19]_0 ),
        .\ex_reg_rs_msb_0_reg[20] (\ex_reg_rs_msb_0_reg[20]_0 ),
        .\ex_reg_rs_msb_0_reg[21] (\ex_reg_rs_msb_0_reg[21]_0 ),
        .\ex_reg_rs_msb_0_reg[22] (\ex_reg_rs_msb_0_reg[22]_0 ),
        .\ex_reg_rs_msb_0_reg[23] (\ex_reg_rs_msb_0_reg[23]_0 ),
        .\ex_reg_rs_msb_0_reg[24] (\ex_reg_rs_msb_0_reg[24]_0 ),
        .\ex_reg_rs_msb_0_reg[25] (\ex_reg_rs_msb_0_reg[25]_0 ),
        .\ex_reg_rs_msb_0_reg[26] (\ex_reg_rs_msb_0_reg[26]_0 ),
        .\ex_reg_rs_msb_0_reg[27] (\ex_reg_rs_msb_0_reg[27]_1 ),
        .\ex_reg_rs_msb_0_reg[8] (\ex_reg_rs_msb_0_reg[8]_0 ),
        .\ex_reg_rs_msb_0_reg[9] (\ex_reg_rs_msb_0_reg[9]_0 ),
        .\ex_reg_rs_msb_1_reg[0] (csr_n_666),
        .\ex_reg_rs_msb_1_reg[1] (csr_n_667),
        .\ex_reg_rs_msb_1_reg[28] (csr_n_678),
        .\ex_reg_rs_msb_1_reg[29] (csr_n_677),
        .\ex_reg_rs_msb_1_reg[2] (csr_n_668),
        .\ex_reg_rs_msb_1_reg[30] (csr_n_676),
        .\ex_reg_rs_msb_1_reg[31] (csr_n_675),
        .\ex_reg_rs_msb_1_reg[32] (csr_n_674),
        .\ex_reg_rs_msb_1_reg[33] (csr_n_673),
        .\ex_reg_rs_msb_1_reg[34] (csr_n_672),
        .\ex_reg_rs_msb_1_reg[35] (csr_n_671),
        .\ex_reg_rs_msb_1_reg[36] (csr_n_670),
        .\ex_reg_rs_msb_1_reg[37] (csr_n_702),
        .\ex_reg_rs_msb_1_reg[38] (csr_n_701),
        .\ex_reg_rs_msb_1_reg[39] (csr_n_700),
        .\ex_reg_rs_msb_1_reg[3] (csr_n_669),
        .\ex_reg_rs_msb_1_reg[40] (csr_n_699),
        .\ex_reg_rs_msb_1_reg[41] (csr_n_698),
        .\ex_reg_rs_msb_1_reg[42] (csr_n_689),
        .\ex_reg_rs_msb_1_reg[43] (csr_n_697),
        .\ex_reg_rs_msb_1_reg[44] (csr_n_696),
        .\ex_reg_rs_msb_1_reg[45] (csr_n_688),
        .\ex_reg_rs_msb_1_reg[46] (csr_n_687),
        .\ex_reg_rs_msb_1_reg[47] (csr_n_686),
        .\ex_reg_rs_msb_1_reg[48] (csr_n_685),
        .\ex_reg_rs_msb_1_reg[49] (csr_n_684),
        .\ex_reg_rs_msb_1_reg[4] (csr_n_642),
        .\ex_reg_rs_msb_1_reg[50] (csr_n_683),
        .\ex_reg_rs_msb_1_reg[51] (csr_n_695),
        .\ex_reg_rs_msb_1_reg[52] (csr_n_694),
        .\ex_reg_rs_msb_1_reg[53] (csr_n_693),
        .\ex_reg_rs_msb_1_reg[54] (csr_n_682),
        .\ex_reg_rs_msb_1_reg[55] (csr_n_681),
        .\ex_reg_rs_msb_1_reg[56] (csr_n_680),
        .\ex_reg_rs_msb_1_reg[57] (csr_n_703),
        .\ex_reg_rs_msb_1_reg[58] (csr_n_692),
        .\ex_reg_rs_msb_1_reg[59] (csr_n_691),
        .\ex_reg_rs_msb_1_reg[5] (csr_n_641),
        .\ex_reg_rs_msb_1_reg[60] (csr_n_690),
        .\ex_reg_rs_msb_1_reg[61] (csr_n_679),
        .\ex_reg_rs_msb_1_reg[6] (csr_n_643),
        .\ex_reg_rs_msb_1_reg[7] (csr_n_644),
        .ex_reg_rvc_reg(ex_reg_rvc_reg_0),
        .ex_reg_valid_reg(ex_reg_valid),
        .ex_reg_xcpt_interrupt0(ex_reg_xcpt_interrupt0),
        .frontend_io_cpu_resp_bits_data(frontend_io_cpu_resp_bits_data),
        .frontend_io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),
        .frontend_io_ptw_pmp_1_cfg_w(frontend_io_ptw_pmp_1_cfg_w),
        .hitsVec_4(hitsVec_4),
        .host_clk(host_clk),
        .ibuf_io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw),
        .ibuf_io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
        .\lrscCount_reg[0] (\lrscCount_reg[0]_0 ),
        .\lrscCount_reg[0]_0 (\lrscCount_reg[0] ),
        .\mem_ctrl_csr_reg[2] (mem_ctrl_csr[2]),
        .mem_ctrl_div(mem_ctrl_div),
        .mem_ctrl_jalr_reg(mem_ctrl_jalr),
        .mem_ctrl_wxd(mem_ctrl_wxd),
        .mem_int_wdata(mem_int_wdata),
        .\mem_reg_cause_reg[1] (mem_reg_cause[1:0]),
        .mem_reg_flush_pipe(mem_reg_flush_pipe),
        .\mem_reg_inst_reg[9] (ibuf_n_52),
        .mem_reg_load(mem_reg_load),
        .mem_reg_sfence_reg(\s1_pc[3]_i_4_n_0 ),
        .mem_reg_sfence_reg_0(\s1_pc[2]_i_4_n_0 ),
        .mem_reg_sfence_reg_1(\s1_pc[4]_i_4_n_0 ),
        .mem_reg_sfence_reg_10(\s1_pc[13]_i_4_n_0 ),
        .mem_reg_sfence_reg_11(\s1_pc[14]_i_4_n_0 ),
        .mem_reg_sfence_reg_12(\s1_pc[15]_i_4_n_0 ),
        .mem_reg_sfence_reg_13(\s1_pc[16]_i_5_n_0 ),
        .mem_reg_sfence_reg_14(\s1_pc[17]_i_4_n_0 ),
        .mem_reg_sfence_reg_15(\s1_pc[18]_i_4_n_0 ),
        .mem_reg_sfence_reg_16(\s1_pc[19]_i_4_n_0 ),
        .mem_reg_sfence_reg_17(\s1_pc[20]_i_5_n_0 ),
        .mem_reg_sfence_reg_18(\s1_pc[21]_i_4_n_0 ),
        .mem_reg_sfence_reg_19(\s1_pc[22]_i_4_n_0 ),
        .mem_reg_sfence_reg_2(\s1_pc[5]_i_3_n_0 ),
        .mem_reg_sfence_reg_20(\s1_pc[23]_i_4_n_0 ),
        .mem_reg_sfence_reg_21(\s1_pc[24]_i_5_n_0 ),
        .mem_reg_sfence_reg_22(\s1_pc[25]_i_4_n_0 ),
        .mem_reg_sfence_reg_23(\s1_pc[26]_i_4_n_0 ),
        .mem_reg_sfence_reg_24(\s1_pc[27]_i_4_n_0 ),
        .mem_reg_sfence_reg_25(\s1_pc[28]_i_5_n_0 ),
        .mem_reg_sfence_reg_26(\s1_pc[29]_i_4_n_0 ),
        .mem_reg_sfence_reg_27(\s1_pc[30]_i_4_n_0 ),
        .mem_reg_sfence_reg_28(\s1_pc[31]_i_4_n_0 ),
        .mem_reg_sfence_reg_29(\s1_pc[32]_i_4_n_0 ),
        .mem_reg_sfence_reg_3(\s1_pc[6]_i_4_n_0 ),
        .mem_reg_sfence_reg_30(\s1_pc[33]_i_3_n_0 ),
        .mem_reg_sfence_reg_31(\s1_pc[34]_i_3_n_0 ),
        .mem_reg_sfence_reg_32(\s1_pc[35]_i_3_n_0 ),
        .mem_reg_sfence_reg_33(\s1_pc[36]_i_4_n_0 ),
        .mem_reg_sfence_reg_34(\s1_pc[37]_i_3_n_0 ),
        .mem_reg_sfence_reg_35(\s1_pc[38]_i_3_n_0 ),
        .mem_reg_sfence_reg_36(\s1_pc[1]_i_3_n_0 ),
        .mem_reg_sfence_reg_37(mem_reg_sfence_reg_2),
        .mem_reg_sfence_reg_38(mem_reg_sfence),
        .mem_reg_sfence_reg_4(\s1_pc[7]_i_4_n_0 ),
        .mem_reg_sfence_reg_5(\s1_pc[8]_i_5_n_0 ),
        .mem_reg_sfence_reg_6(\s1_pc[9]_i_4_n_0 ),
        .mem_reg_sfence_reg_7(\s1_pc[10]_i_4_n_0 ),
        .mem_reg_sfence_reg_8(\s1_pc[11]_i_4_n_0 ),
        .mem_reg_sfence_reg_9(\s1_pc[12]_i_5_n_0 ),
        .mem_reg_slow_bypass_reg(ibuf_n_68),
        .mem_reg_store(mem_reg_store),
        .mem_reg_valid_reg(mem_reg_replay_reg_0),
        .mem_reg_valid_reg_0(mem_reg_valid),
        .mem_reg_xcpt_interrupt_reg(mem_reg_xcpt_interrupt),
        .mem_reg_xcpt_reg(mem_reg_xcpt),
        .nBufValid_reg(nBufValid_reg_0),
        .nBufValid_reg_0(nBufValid_reg_1),
        .nBufValid_reg_1(\ex_ctrl_sel_alu2_reg[1]_3 ),
        .nBufValid_reg_2(ibuf_n_47),
        .nBufValid_reg_3(nBufValid_reg_2),
        .p_0_in(p_0_in),
        .p_13_in(p_13_in),
        .q_reg(q_reg),
        .\r_pte_ppn_reg[0] (\r_pte_ppn_reg[0] ),
        .\r_pte_ppn_reg[10] (\r_pte_ppn_reg[10] ),
        .\r_pte_ppn_reg[11] (\r_pte_ppn_reg[11] ),
        .\r_pte_ppn_reg[12] (\r_pte_ppn_reg[12] ),
        .\r_pte_ppn_reg[13] (\r_pte_ppn_reg[13] ),
        .\r_pte_ppn_reg[14] (\r_pte_ppn_reg[14] ),
        .\r_pte_ppn_reg[15] (\r_pte_ppn_reg[15] ),
        .\r_pte_ppn_reg[16] (\r_pte_ppn_reg[16] ),
        .\r_pte_ppn_reg[16]_0 (\r_pte_ppn_reg[16]_0 ),
        .\r_pte_ppn_reg[16]_1 (\r_pte_ppn_reg[16]_1 ),
        .\r_pte_ppn_reg[16]_2 (\r_pte_ppn_reg[16]_2 ),
        .\r_pte_ppn_reg[16]_3 (\r_pte_ppn_reg[16]_3 ),
        .\r_pte_ppn_reg[16]_4 (\r_pte_ppn_reg[16]_4 ),
        .\r_pte_ppn_reg[16]_5 (\r_pte_ppn_reg[16]_5 ),
        .\r_pte_ppn_reg[16]_6 (\r_pte_ppn_reg[16]_6 ),
        .\r_pte_ppn_reg[16]_7 (\r_pte_ppn_reg[16]_7 ),
        .\r_pte_ppn_reg[17] (\r_pte_ppn_reg[17] ),
        .\r_pte_ppn_reg[18] (\r_pte_ppn_reg[18] ),
        .\r_pte_ppn_reg[19] (\r_pte_ppn_reg[19] ),
        .\r_pte_ppn_reg[19]_0 (\r_pte_ppn_reg[19]_0 ),
        .\r_pte_ppn_reg[1] (\r_pte_ppn_reg[1] ),
        .\r_pte_ppn_reg[2] (\r_pte_ppn_reg[2] ),
        .\r_pte_ppn_reg[3] (\r_pte_ppn_reg[3] ),
        .\r_pte_ppn_reg[3]_0 (\r_pte_ppn_reg[3]_0 ),
        .\r_pte_ppn_reg[3]_1 (\r_pte_ppn_reg[3]_1 ),
        .\r_pte_ppn_reg[3]_2 (\r_pte_ppn_reg[3]_2 ),
        .\r_pte_ppn_reg[3]_3 (\r_pte_ppn_reg[3]_3 ),
        .\r_pte_ppn_reg[3]_4 (\r_pte_ppn_reg[3]_4 ),
        .\r_pte_ppn_reg[3]_5 (\r_pte_ppn_reg[3]_5 ),
        .\r_pte_ppn_reg[3]_6 (\r_pte_ppn_reg[3]_6 ),
        .\r_pte_ppn_reg[3]_7 (\r_pte_ppn_reg[3]_7 ),
        .\r_pte_ppn_reg[4] (\r_pte_ppn_reg[4] ),
        .\r_pte_ppn_reg[5] (\r_pte_ppn_reg[5] ),
        .\r_pte_ppn_reg[5]_0 (\r_pte_ppn_reg[5]_0 ),
        .\r_pte_ppn_reg[5]_1 (\r_pte_ppn_reg[5]_1 ),
        .\r_pte_ppn_reg[5]_2 (\r_pte_ppn_reg[5]_2 ),
        .\r_pte_ppn_reg[5]_3 (\r_pte_ppn_reg[5]_3 ),
        .\r_pte_ppn_reg[5]_4 (\r_pte_ppn_reg[5]_4 ),
        .\r_pte_ppn_reg[5]_5 (\r_pte_ppn_reg[5]_5 ),
        .\r_pte_ppn_reg[5]_6 (\r_pte_ppn_reg[5]_6 ),
        .\r_pte_ppn_reg[5]_7 (\r_pte_ppn_reg[5]_7 ),
        .\r_pte_ppn_reg[6] (\r_pte_ppn_reg[6] ),
        .\r_pte_ppn_reg[7] (\r_pte_ppn_reg[7] ),
        .\r_pte_ppn_reg[7]_0 (\r_pte_ppn_reg[7]_0 ),
        .\r_pte_ppn_reg[7]_1 (\r_pte_ppn_reg[7]_1 ),
        .\r_pte_ppn_reg[7]_2 (\r_pte_ppn_reg[7]_2 ),
        .\r_pte_ppn_reg[7]_3 (\r_pte_ppn_reg[7]_3 ),
        .\r_pte_ppn_reg[7]_4 (\r_pte_ppn_reg[7]_4 ),
        .\r_pte_ppn_reg[7]_5 (\r_pte_ppn_reg[7]_5 ),
        .\r_pte_ppn_reg[7]_6 (\r_pte_ppn_reg[7]_6 ),
        .\r_pte_ppn_reg[7]_7 (\r_pte_ppn_reg[7]_7 ),
        .\r_pte_ppn_reg[8] (\r_pte_ppn_reg[8] ),
        .\r_pte_ppn_reg[9] (\r_pte_ppn_reg[9] ),
        .\r_refill_waddr_reg[0] (\r_refill_waddr_reg[0] ),
        .\r_refill_waddr_reg[1] (\r_refill_waddr_reg[1] ),
        .\reg_bp_0_address_reg[36]_0 (\reg_bp_0_address_reg[36] ),
        .\reg_bp_0_address_reg[3]_0 (\reg_bp_0_address_reg[3] ),
        .reg_bp_0_control_action_reg_0(reg_bp_0_control_action_reg),
        .reg_bp_0_control_action_reg_1(ibuf_n_65),
        .\reg_bp_0_control_tmatch_reg[1]_0 (\reg_bp_0_control_tmatch_reg[1]_0 ),
        .\reg_dcsr_cause_reg[0]_0 (\reg_dcsr_cause_reg[0] ),
        .\reg_dcsr_cause_reg[1]_0 (\reg_dcsr_cause_reg[1] ),
        .reg_debug_reg_0(reg_dcsr_prv),
        .reg_debug_reg_1(reg_debug_reg_0),
        .reg_debug_reg_2(reg_debug_reg_1),
        .reg_debug_reg_3(reg_debug_reg_2),
        .\reg_dpc_reg[12]_0 (\reg_dpc_reg[12] ),
        .\reg_dscratch_reg[0]_0 (\reg_dscratch_reg[0] ),
        .\reg_entries_0_reg[0] (\reg_entries_0_reg[0] ),
        .\reg_entries_0_reg[0]_0 (\reg_entries_0_reg[0]_0 ),
        .\reg_entries_0_reg[0]_1 (\reg_entries_0_reg[0]_1 ),
        .\reg_entries_0_reg[0]_2 (\reg_entries_0_reg[0]_2 ),
        .\reg_entries_0_reg[0]_3 (\reg_entries_0_reg[0]_3 ),
        .\reg_entries_0_reg[0]_4 (\reg_entries_0_reg[0]_4 ),
        .\reg_entries_0_reg[0]_5 (\reg_entries_0_reg[0]_5 ),
        .\reg_entries_0_reg[0]_6 (\reg_entries_0_reg[0]_6 ),
        .\reg_entries_0_reg[0]_7 (\reg_entries_0_reg[0]_7 ),
        .\reg_entries_0_reg[10] (\reg_entries_0_reg[10] ),
        .\reg_entries_0_reg[4] (\reg_entries_0_reg[4] ),
        .\reg_entries_0_reg[4]_0 (\reg_entries_0_reg[4]_0 ),
        .\reg_entries_0_reg[4]_1 (\reg_entries_0_reg[4]_1 ),
        .\reg_entries_0_reg[4]_10 (\reg_entries_0_reg[4]_10 ),
        .\reg_entries_0_reg[4]_11 (\reg_entries_0_reg[4]_11 ),
        .\reg_entries_0_reg[4]_12 (\reg_entries_0_reg[4]_12 ),
        .\reg_entries_0_reg[4]_13 (\reg_entries_0_reg[4]_13 ),
        .\reg_entries_0_reg[4]_14 (\reg_entries_0_reg[4]_14 ),
        .\reg_entries_0_reg[4]_15 (\reg_entries_0_reg[4]_15 ),
        .\reg_entries_0_reg[4]_16 (\reg_entries_0_reg[4]_16 ),
        .\reg_entries_0_reg[4]_17 (\reg_entries_0_reg[4]_17 ),
        .\reg_entries_0_reg[4]_18 (\reg_entries_0_reg[4]_18 ),
        .\reg_entries_0_reg[4]_19 (\reg_entries_0_reg[4]_19 ),
        .\reg_entries_0_reg[4]_2 (\reg_entries_0_reg[4]_2 ),
        .\reg_entries_0_reg[4]_20 (\reg_entries_0_reg[4]_20 ),
        .\reg_entries_0_reg[4]_21 (\reg_entries_0_reg[4]_21 ),
        .\reg_entries_0_reg[4]_22 (\reg_entries_0_reg[4]_22 ),
        .\reg_entries_0_reg[4]_23 (\reg_entries_0_reg[4]_23 ),
        .\reg_entries_0_reg[4]_24 (\reg_entries_0_reg[4]_24 ),
        .\reg_entries_0_reg[4]_25 (\reg_entries_0_reg[4]_25 ),
        .\reg_entries_0_reg[4]_3 (\reg_entries_0_reg[4]_3 ),
        .\reg_entries_0_reg[4]_4 (\reg_entries_0_reg[4]_4 ),
        .\reg_entries_0_reg[4]_5 (\reg_entries_0_reg[4]_5 ),
        .\reg_entries_0_reg[4]_6 (\reg_entries_0_reg[4]_6 ),
        .\reg_entries_0_reg[4]_7 (\reg_entries_0_reg[4]_7 ),
        .\reg_entries_0_reg[4]_8 (\reg_entries_0_reg[4]_8 ),
        .\reg_entries_0_reg[4]_9 (\reg_entries_0_reg[4]_9 ),
        .\reg_entries_0_reg[5] (\reg_entries_0_reg[5] ),
        .\reg_entries_0_reg[5]_0 (\reg_entries_0_reg[5]_0 ),
        .\reg_entries_0_reg[5]_1 (\reg_entries_0_reg[5]_1 ),
        .\reg_entries_0_reg[5]_10 (\reg_entries_0_reg[5]_10 ),
        .\reg_entries_0_reg[5]_11 (\reg_entries_0_reg[5]_11 ),
        .\reg_entries_0_reg[5]_12 (\reg_entries_0_reg[5]_12 ),
        .\reg_entries_0_reg[5]_13 (\reg_entries_0_reg[5]_13 ),
        .\reg_entries_0_reg[5]_14 (\reg_entries_0_reg[5]_14 ),
        .\reg_entries_0_reg[5]_15 (\reg_entries_0_reg[5]_15 ),
        .\reg_entries_0_reg[5]_16 (\reg_entries_0_reg[5]_16 ),
        .\reg_entries_0_reg[5]_17 (\reg_entries_0_reg[5]_17 ),
        .\reg_entries_0_reg[5]_18 (\reg_entries_0_reg[5]_18 ),
        .\reg_entries_0_reg[5]_19 (\reg_entries_0_reg[5]_19 ),
        .\reg_entries_0_reg[5]_2 (\reg_entries_0_reg[5]_2 ),
        .\reg_entries_0_reg[5]_20 (\reg_entries_0_reg[5]_20 ),
        .\reg_entries_0_reg[5]_21 (\reg_entries_0_reg[5]_21 ),
        .\reg_entries_0_reg[5]_22 (\reg_entries_0_reg[5]_22 ),
        .\reg_entries_0_reg[5]_23 (\reg_entries_0_reg[5]_23 ),
        .\reg_entries_0_reg[5]_24 (\reg_entries_0_reg[5]_24 ),
        .\reg_entries_0_reg[5]_25 (\reg_entries_0_reg[5]_25 ),
        .\reg_entries_0_reg[5]_26 (\reg_entries_0_reg[5]_26 ),
        .\reg_entries_0_reg[5]_27 (\reg_entries_0_reg[5]_27 ),
        .\reg_entries_0_reg[5]_28 (\reg_entries_0_reg[5]_28 ),
        .\reg_entries_0_reg[5]_29 (\reg_entries_0_reg[5]_29 ),
        .\reg_entries_0_reg[5]_3 (\reg_entries_0_reg[5]_3 ),
        .\reg_entries_0_reg[5]_30 (\reg_entries_0_reg[5]_30 ),
        .\reg_entries_0_reg[5]_31 (\reg_entries_0_reg[5]_31 ),
        .\reg_entries_0_reg[5]_32 (\reg_entries_0_reg[5]_32 ),
        .\reg_entries_0_reg[5]_33 (\reg_entries_0_reg[5]_33 ),
        .\reg_entries_0_reg[5]_34 (\reg_entries_0_reg[5]_34 ),
        .\reg_entries_0_reg[5]_35 (\reg_entries_0_reg[5]_35 ),
        .\reg_entries_0_reg[5]_36 (\reg_entries_0_reg[5]_36 ),
        .\reg_entries_0_reg[5]_37 (\reg_entries_0_reg[5]_37 ),
        .\reg_entries_0_reg[5]_38 (\reg_entries_0_reg[5]_38 ),
        .\reg_entries_0_reg[5]_39 (\reg_entries_0_reg[5]_39 ),
        .\reg_entries_0_reg[5]_4 (\reg_entries_0_reg[5]_4 ),
        .\reg_entries_0_reg[5]_40 (\reg_entries_0_reg[5]_40 ),
        .\reg_entries_0_reg[5]_41 (\reg_entries_0_reg[5]_41 ),
        .\reg_entries_0_reg[5]_42 (\reg_entries_0_reg[5]_42 ),
        .\reg_entries_0_reg[5]_43 (\reg_entries_0_reg[5]_43 ),
        .\reg_entries_0_reg[5]_44 (\reg_entries_0_reg[5]_44 ),
        .\reg_entries_0_reg[5]_45 (\reg_entries_0_reg[5]_45 ),
        .\reg_entries_0_reg[5]_46 (\reg_entries_0_reg[5]_46 ),
        .\reg_entries_0_reg[5]_47 (\reg_entries_0_reg[5]_47 ),
        .\reg_entries_0_reg[5]_5 (\reg_entries_0_reg[5]_5 ),
        .\reg_entries_0_reg[5]_6 (\reg_entries_0_reg[5]_6 ),
        .\reg_entries_0_reg[5]_7 (\reg_entries_0_reg[5]_7 ),
        .\reg_entries_0_reg[5]_8 (\reg_entries_0_reg[5]_8 ),
        .\reg_entries_0_reg[5]_9 (\reg_entries_0_reg[5]_9 ),
        .\reg_entries_0_reg[6] (\reg_entries_0_reg[6] ),
        .\reg_entries_0_reg[6]_0 (\reg_entries_0_reg[6]_0 ),
        .\reg_entries_0_reg[6]_1 (\reg_entries_0_reg[6]_1 ),
        .\reg_entries_0_reg[6]_10 (\reg_entries_0_reg[6]_10 ),
        .\reg_entries_0_reg[6]_11 (\reg_entries_0_reg[6]_11 ),
        .\reg_entries_0_reg[6]_12 (\reg_entries_0_reg[6]_12 ),
        .\reg_entries_0_reg[6]_13 (\reg_entries_0_reg[6]_13 ),
        .\reg_entries_0_reg[6]_14 (\reg_entries_0_reg[6]_14 ),
        .\reg_entries_0_reg[6]_15 (\reg_entries_0_reg[6]_15 ),
        .\reg_entries_0_reg[6]_16 (\reg_entries_0_reg[6]_16 ),
        .\reg_entries_0_reg[6]_17 (\reg_entries_0_reg[6]_17 ),
        .\reg_entries_0_reg[6]_18 (\reg_entries_0_reg[6]_18 ),
        .\reg_entries_0_reg[6]_19 (\reg_entries_0_reg[6]_19 ),
        .\reg_entries_0_reg[6]_2 (\reg_entries_0_reg[6]_2 ),
        .\reg_entries_0_reg[6]_20 (\reg_entries_0_reg[6]_20 ),
        .\reg_entries_0_reg[6]_21 (\reg_entries_0_reg[6]_21 ),
        .\reg_entries_0_reg[6]_22 (\reg_entries_0_reg[6]_22 ),
        .\reg_entries_0_reg[6]_23 (\reg_entries_0_reg[6]_23 ),
        .\reg_entries_0_reg[6]_24 (\reg_entries_0_reg[6]_24 ),
        .\reg_entries_0_reg[6]_25 (\reg_entries_0_reg[6]_25 ),
        .\reg_entries_0_reg[6]_26 (\reg_entries_0_reg[6]_26 ),
        .\reg_entries_0_reg[6]_27 (\reg_entries_0_reg[6]_27 ),
        .\reg_entries_0_reg[6]_28 (\reg_entries_0_reg[6]_28 ),
        .\reg_entries_0_reg[6]_29 (\reg_entries_0_reg[6]_29 ),
        .\reg_entries_0_reg[6]_3 (\reg_entries_0_reg[6]_3 ),
        .\reg_entries_0_reg[6]_30 (\reg_entries_0_reg[6]_30 ),
        .\reg_entries_0_reg[6]_31 (\reg_entries_0_reg[6]_31 ),
        .\reg_entries_0_reg[6]_32 (\reg_entries_0_reg[6]_32 ),
        .\reg_entries_0_reg[6]_33 (\reg_entries_0_reg[6]_33 ),
        .\reg_entries_0_reg[6]_34 (\reg_entries_0_reg[6]_34 ),
        .\reg_entries_0_reg[6]_35 (\reg_entries_0_reg[6]_35 ),
        .\reg_entries_0_reg[6]_36 (\reg_entries_0_reg[6]_36 ),
        .\reg_entries_0_reg[6]_37 (\reg_entries_0_reg[6]_37 ),
        .\reg_entries_0_reg[6]_38 (\reg_entries_0_reg[6]_38 ),
        .\reg_entries_0_reg[6]_39 (\reg_entries_0_reg[6]_39 ),
        .\reg_entries_0_reg[6]_4 (\reg_entries_0_reg[6]_4 ),
        .\reg_entries_0_reg[6]_40 (\reg_entries_0_reg[6]_40 ),
        .\reg_entries_0_reg[6]_41 (\reg_entries_0_reg[6]_41 ),
        .\reg_entries_0_reg[6]_42 (\reg_entries_0_reg[6]_42 ),
        .\reg_entries_0_reg[6]_43 (\reg_entries_0_reg[6]_43 ),
        .\reg_entries_0_reg[6]_44 (\reg_entries_0_reg[6]_44 ),
        .\reg_entries_0_reg[6]_45 (\reg_entries_0_reg[6]_45 ),
        .\reg_entries_0_reg[6]_46 (\reg_entries_0_reg[6]_46 ),
        .\reg_entries_0_reg[6]_47 (\reg_entries_0_reg[6]_47 ),
        .\reg_entries_0_reg[6]_48 (\reg_entries_0_reg[6]_48 ),
        .\reg_entries_0_reg[6]_49 (\reg_entries_0_reg[6]_49 ),
        .\reg_entries_0_reg[6]_5 (\reg_entries_0_reg[6]_5 ),
        .\reg_entries_0_reg[6]_50 (\reg_entries_0_reg[6]_50 ),
        .\reg_entries_0_reg[6]_51 (\reg_entries_0_reg[6]_51 ),
        .\reg_entries_0_reg[6]_52 (\reg_entries_0_reg[6]_52 ),
        .\reg_entries_0_reg[6]_53 (\reg_entries_0_reg[6]_53 ),
        .\reg_entries_0_reg[6]_54 (\reg_entries_0_reg[6]_54 ),
        .\reg_entries_0_reg[6]_55 (\reg_entries_0_reg[6]_55 ),
        .\reg_entries_0_reg[6]_56 (\reg_entries_0_reg[6]_56 ),
        .\reg_entries_0_reg[6]_57 (\reg_entries_0_reg[6]_57 ),
        .\reg_entries_0_reg[6]_6 (\reg_entries_0_reg[6]_6 ),
        .\reg_entries_0_reg[6]_7 (\reg_entries_0_reg[6]_7 ),
        .\reg_entries_0_reg[6]_8 (\reg_entries_0_reg[6]_8 ),
        .\reg_entries_0_reg[6]_9 (\reg_entries_0_reg[6]_9 ),
        .\reg_entries_1_reg[0] (\reg_entries_1_reg[0] ),
        .\reg_entries_1_reg[0]_0 (\reg_entries_1_reg[0]_0 ),
        .\reg_entries_1_reg[0]_1 (\reg_entries_1_reg[0]_1 ),
        .\reg_entries_1_reg[0]_10 (\reg_entries_1_reg[0]_11 ),
        .\reg_entries_1_reg[0]_11 (\reg_entries_1_reg[0]_12 ),
        .\reg_entries_1_reg[0]_12 (\reg_entries_1_reg[0]_13 ),
        .\reg_entries_1_reg[0]_13 (\reg_entries_1_reg[0]_8 ),
        .\reg_entries_1_reg[0]_14 (\reg_entries_1_reg[0]_14 ),
        .\reg_entries_1_reg[0]_15 (\reg_entries_1_reg[0]_15 ),
        .\reg_entries_1_reg[0]_16 (\reg_entries_1_reg[0]_16 ),
        .\reg_entries_1_reg[0]_17 (\reg_entries_1_reg[0]_17 ),
        .\reg_entries_1_reg[0]_18 (\reg_entries_1_reg[0]_18 ),
        .\reg_entries_1_reg[0]_19 (\reg_entries_1_reg[0]_19 ),
        .\reg_entries_1_reg[0]_2 (\reg_entries_1_reg[0]_2 ),
        .\reg_entries_1_reg[0]_20 (\reg_entries_1_reg[0]_20 ),
        .\reg_entries_1_reg[0]_21 (\reg_entries_1_reg[0]_21 ),
        .\reg_entries_1_reg[0]_22 (\reg_entries_1_reg[0]_22 ),
        .\reg_entries_1_reg[0]_23 (\reg_entries_1_reg[0]_23 ),
        .\reg_entries_1_reg[0]_24 (\reg_entries_1_reg[0]_24 ),
        .\reg_entries_1_reg[0]_25 (\reg_entries_1_reg[0]_25 ),
        .\reg_entries_1_reg[0]_26 (\reg_entries_1_reg[0]_26 ),
        .\reg_entries_1_reg[0]_27 (\reg_entries_1_reg[0]_27 ),
        .\reg_entries_1_reg[0]_28 (\reg_entries_1_reg[0]_28 ),
        .\reg_entries_1_reg[0]_29 (\reg_entries_1_reg[0]_29 ),
        .\reg_entries_1_reg[0]_3 (\reg_entries_1_reg[0]_3 ),
        .\reg_entries_1_reg[0]_30 (\reg_entries_1_reg[0]_30 ),
        .\reg_entries_1_reg[0]_31 (\reg_entries_1_reg[0]_31 ),
        .\reg_entries_1_reg[0]_32 (\reg_entries_1_reg[0]_32 ),
        .\reg_entries_1_reg[0]_33 (\reg_entries_1_reg[0]_33 ),
        .\reg_entries_1_reg[0]_34 (\reg_entries_1_reg[0]_34 ),
        .\reg_entries_1_reg[0]_35 (\reg_entries_1_reg[0]_35 ),
        .\reg_entries_1_reg[0]_36 (\reg_entries_1_reg[0]_36 ),
        .\reg_entries_1_reg[0]_37 (\reg_entries_1_reg[0]_37 ),
        .\reg_entries_1_reg[0]_38 (\reg_entries_1_reg[0]_38 ),
        .\reg_entries_1_reg[0]_39 (\reg_entries_1_reg[0]_39 ),
        .\reg_entries_1_reg[0]_4 (\reg_entries_1_reg[0]_4 ),
        .\reg_entries_1_reg[0]_40 (\reg_entries_1_reg[0]_40 ),
        .\reg_entries_1_reg[0]_41 (\reg_entries_1_reg[0]_41 ),
        .\reg_entries_1_reg[0]_42 (\reg_entries_1_reg[0]_42 ),
        .\reg_entries_1_reg[0]_43 (\reg_entries_1_reg[0]_43 ),
        .\reg_entries_1_reg[0]_44 (\reg_entries_1_reg[0]_44 ),
        .\reg_entries_1_reg[0]_45 (\reg_entries_1_reg[0]_45 ),
        .\reg_entries_1_reg[0]_46 (\reg_entries_1_reg[0]_46 ),
        .\reg_entries_1_reg[0]_47 (\reg_entries_1_reg[0]_47 ),
        .\reg_entries_1_reg[0]_5 (\reg_entries_1_reg[0]_5 ),
        .\reg_entries_1_reg[0]_6 (\reg_entries_1_reg[0]_6 ),
        .\reg_entries_1_reg[0]_7 (\reg_entries_1_reg[0]_7 ),
        .\reg_entries_1_reg[0]_8 (\reg_entries_1_reg[0]_9 ),
        .\reg_entries_1_reg[0]_9 (\reg_entries_1_reg[0]_10 ),
        .\reg_entries_1_reg[12] (\reg_entries_1_reg[12] ),
        .\reg_entries_2_reg[12] (\reg_entries_2_reg[12] ),
        .\reg_entries_3_reg[11] (\reg_entries_3_reg[11] ),
        .\reg_entries_3_reg[12] (\reg_entries_3_reg[12] ),
        .\reg_entries_4_reg[61] (\reg_entries_4_reg[61] ),
        .\reg_entries_4_reg[61]_0 (\reg_entries_4_reg[61]_0 ),
        .\reg_mbadaddr_reg[12]_0 (\reg_mbadaddr_reg[12] ),
        .\reg_mcause_reg[0]_0 (\reg_mcause_reg[0] ),
        .\reg_mepc_reg[12]_0 (\reg_mepc_reg[12] ),
        .\reg_mie_reg[7]_0 (\reg_mie_reg[7] ),
        .reg_mip_seip_reg_0(reg_mip_seip_reg),
        .\reg_misa_reg[0]_0 (\reg_misa_reg[0] ),
        .\reg_misa_reg[12]_0 (\reg_misa_reg[12] [1]),
        .reg_mstatus_mie(reg_mstatus_mie),
        .reg_mstatus_mie_reg_0(reg_mstatus_mie_reg),
        .reg_mstatus_mie_reg_1(reg_mstatus_mie_reg_0),
        .reg_mstatus_mpie_reg_0(reg_mstatus_mpie_reg),
        .reg_mstatus_mpie_reg_1(reg_mstatus_mpie_reg_0),
        .\reg_mstatus_mpp_reg[0]_0 (\reg_mstatus_mpp_reg[0] ),
        .\reg_mstatus_mpp_reg[1]_0 (\reg_mstatus_mpp_reg[1] ),
        .reg_mstatus_mxr_reg_0(dcache_io_ptw_status_mxr),
        .\reg_mstatus_prv_reg[0]_0 (frontend_io_ptw_status_prv[0]),
        .\reg_mstatus_prv_reg[1]_0 (frontend_io_ptw_status_prv[1]),
        .\reg_mstatus_prv_reg[1]_1 (\reg_mstatus_prv_reg[1] ),
        .\reg_mstatus_prv_reg[1]_2 (\reg_mstatus_prv_reg[1]_0 ),
        .\reg_mstatus_prv_reg[1]_3 (\reg_mstatus_prv_reg[1]_1 ),
        .\reg_mstatus_prv_reg[1]_4 (\reg_mstatus_prv_reg[1]_2 ),
        .reg_mstatus_spie_reg_0(reg_mstatus_spie_reg),
        .reg_mstatus_sum_reg_0(dcache_io_ptw_status_sum),
        .\reg_mtvec_reg[20]_0 (\reg_mtvec_reg[20] ),
        .\reg_mtvec_reg[21]_0 (\reg_mtvec_reg[21] ),
        .\reg_mtvec_reg[22]_0 (\reg_mtvec_reg[22] ),
        .\reg_mtvec_reg[29]_0 (\reg_mtvec_reg[29]_0 ),
        .\reg_mtvec_reg[29]_1 (\reg_mtvec_reg[29]_1 ),
        .\reg_mtvec_reg[29]_2 (\reg_mtvec_reg[29]_2 ),
        .\reg_mtvec_reg[29]_3 (\reg_mtvec_reg[29]_3 ),
        .\reg_mtvec_reg[29]_4 (\reg_mtvec_reg[29]_4 ),
        .\reg_mtvec_reg[29]_5 (\reg_mtvec_reg[29]_5 ),
        .\reg_mtvec_reg[29]_6 (\reg_mtvec_reg[29]_6 ),
        .\reg_mtvec_reg[4]_0 (\reg_mtvec_reg[4] ),
        .\reg_pmp_0_addr_reg[13]_0 (\reg_pmp_0_addr_reg[13] ),
        .\reg_pmp_0_addr_reg[17]_0 (\reg_pmp_0_addr_reg[17] ),
        .\reg_pmp_0_addr_reg[19]_0 (\reg_pmp_0_addr_reg[19] ),
        .\reg_pmp_0_addr_reg[23]_0 (\reg_pmp_0_addr_reg[23] ),
        .\reg_pmp_0_addr_reg[28]_0 (\reg_pmp_0_addr_reg[28] ),
        .\reg_pmp_0_addr_reg[28]_1 (\reg_pmp_0_addr_reg[28]_0 ),
        .\reg_pmp_0_addr_reg[29]_0 (\reg_pmp_0_addr_reg[29] ),
        .\reg_pmp_0_addr_reg[29]_1 (\reg_pmp_0_addr_reg[29]_0 ),
        .\reg_pmp_1_addr_reg[13]_0 (\reg_pmp_1_addr_reg[13] ),
        .\reg_pmp_1_addr_reg[17]_0 (\reg_pmp_1_addr_reg[17] ),
        .\reg_pmp_1_addr_reg[19]_0 (\reg_pmp_1_addr_reg[19] ),
        .\reg_pmp_1_addr_reg[28]_0 (\reg_pmp_1_addr_reg[28] ),
        .\reg_pmp_1_addr_reg[28]_1 (\reg_pmp_1_addr_reg[28]_0 ),
        .\reg_pmp_1_addr_reg[29]_0 (\reg_pmp_1_addr_reg[29] ),
        .\reg_pmp_1_addr_reg[29]_1 (\reg_pmp_1_addr_reg[29]_0 ),
        .\reg_pmp_1_cfg_a_reg[0]_0 (frontend_io_ptw_pmp_1_cfg_a[0]),
        .\reg_pmp_1_cfg_a_reg[0]_1 (\reg_pmp_1_cfg_a_reg[0] ),
        .\reg_pmp_1_cfg_a_reg[1]_0 (frontend_io_ptw_pmp_1_cfg_a[1]),
        .reg_pmp_1_cfg_w_reg_0(reg_pmp_1_cfg_w_reg),
        .\reg_pmp_2_addr_reg[0]_0 (\reg_pmp_2_addr_reg[0] ),
        .\reg_pmp_2_addr_reg[13]_0 (\reg_pmp_2_addr_reg[13] ),
        .\reg_pmp_2_addr_reg[17]_0 (\reg_pmp_2_addr_reg[17] ),
        .\reg_pmp_2_addr_reg[19]_0 (\reg_pmp_2_addr_reg[19] ),
        .\reg_pmp_2_addr_reg[28]_0 (\reg_pmp_2_addr_reg[28] ),
        .\reg_pmp_2_addr_reg[28]_1 (\reg_pmp_2_addr_reg[28]_0 ),
        .\reg_pmp_2_addr_reg[29]_0 (\reg_pmp_2_addr_reg[29] ),
        .\reg_pmp_2_addr_reg[29]_1 (\reg_pmp_2_addr_reg[29]_0 ),
        .\reg_pmp_2_addr_reg[29]_2 (\reg_pmp_2_addr_reg[29]_1 ),
        .\reg_pmp_2_cfg_a_reg[0]_0 (frontend_io_ptw_pmp_2_cfg_a[0]),
        .\reg_pmp_2_cfg_a_reg[0]_1 (\reg_pmp_2_cfg_a_reg[0] ),
        .\reg_pmp_2_cfg_a_reg[1]_0 (frontend_io_ptw_pmp_2_cfg_a[1]),
        .\reg_pmp_3_addr_reg[13]_0 (\reg_pmp_3_addr_reg[13] ),
        .\reg_pmp_3_addr_reg[17]_0 (\reg_pmp_3_addr_reg[17] ),
        .\reg_pmp_3_addr_reg[18]_0 (\reg_pmp_3_addr_reg[18] ),
        .\reg_pmp_3_addr_reg[19]_0 (\reg_pmp_3_addr_reg[19] ),
        .\reg_pmp_3_addr_reg[23]_0 (\reg_pmp_3_addr_reg[23] ),
        .\reg_pmp_3_addr_reg[28]_0 (\reg_pmp_3_addr_reg[28] ),
        .\reg_pmp_3_addr_reg[28]_1 (\reg_pmp_3_addr_reg[28]_0 ),
        .\reg_pmp_3_addr_reg[29]_0 (\reg_pmp_3_addr_reg[29] ),
        .\reg_pmp_3_addr_reg[29]_1 (\reg_pmp_3_addr_reg[29]_0 ),
        .\reg_pmp_3_addr_reg[29]_2 (\reg_pmp_3_addr_reg[29]_1 ),
        .\reg_pmp_4_addr_reg[0]_0 (\reg_pmp_4_addr_reg[0] ),
        .\reg_pmp_4_addr_reg[13]_0 (\reg_pmp_4_addr_reg[13] ),
        .\reg_pmp_4_addr_reg[14]_0 (\reg_pmp_4_addr_reg[14] ),
        .\reg_pmp_4_addr_reg[17]_0 (\reg_pmp_4_addr_reg[17] ),
        .\reg_pmp_4_addr_reg[19]_0 (\reg_pmp_4_addr_reg[19] ),
        .\reg_pmp_4_addr_reg[28]_0 (\reg_pmp_4_addr_reg[28] ),
        .\reg_pmp_4_addr_reg[28]_1 (\reg_pmp_4_addr_reg[28]_0 ),
        .\reg_pmp_4_addr_reg[29]_0 (\reg_pmp_4_addr_reg[29] ),
        .\reg_pmp_4_addr_reg[29]_1 (\reg_pmp_4_addr_reg[29]_0 ),
        .\reg_pmp_4_cfg_a_reg[1]_0 (\reg_pmp_4_cfg_a_reg[1] ),
        .\reg_pmp_5_addr_reg[13]_0 (\reg_pmp_5_addr_reg[13] ),
        .\reg_pmp_5_addr_reg[17]_0 (\reg_pmp_5_addr_reg[17] ),
        .\reg_pmp_5_addr_reg[19]_0 (\reg_pmp_5_addr_reg[19] ),
        .\reg_pmp_5_addr_reg[20]_0 (\reg_pmp_5_addr_reg[20] ),
        .\reg_pmp_5_addr_reg[28]_0 (\reg_pmp_5_addr_reg[28] ),
        .\reg_pmp_5_addr_reg[28]_1 (\reg_pmp_5_addr_reg[28]_0 ),
        .\reg_pmp_5_addr_reg[29]_0 (\reg_pmp_5_addr_reg[29] ),
        .\reg_pmp_5_addr_reg[29]_1 (\reg_pmp_5_addr_reg[29]_0 ),
        .\reg_pmp_5_cfg_a_reg[1]_0 (\reg_pmp_5_cfg_a_reg[1] ),
        .\reg_pmp_5_cfg_a_reg[1]_1 (\reg_pmp_5_cfg_a_reg[1]_0 ),
        .\reg_pmp_6_addr_reg[13]_0 (\reg_pmp_6_addr_reg[13] ),
        .\reg_pmp_6_addr_reg[17]_0 (\reg_pmp_6_addr_reg[17] ),
        .\reg_pmp_6_addr_reg[19]_0 (\reg_pmp_6_addr_reg[19] ),
        .\reg_pmp_6_addr_reg[28]_0 (\reg_pmp_6_addr_reg[28] ),
        .\reg_pmp_6_addr_reg[28]_1 (\reg_pmp_6_addr_reg[28]_0 ),
        .\reg_pmp_6_addr_reg[29]_0 (\reg_pmp_6_addr_reg[29] ),
        .\reg_pmp_6_addr_reg[29]_1 (\reg_pmp_6_addr_reg[29]_0 ),
        .\reg_pmp_6_cfg_a_reg[0]_0 (frontend_io_ptw_pmp_6_cfg_a[0]),
        .\reg_pmp_6_cfg_a_reg[1]_0 (frontend_io_ptw_pmp_6_cfg_a[1]),
        .\reg_pmp_7_addr_reg[13]_0 (\reg_pmp_7_addr_reg[13] ),
        .\reg_pmp_7_addr_reg[17]_0 (\reg_pmp_7_addr_reg[17] ),
        .\reg_pmp_7_addr_reg[17]_1 (\reg_pmp_7_addr_reg[17]_0 ),
        .\reg_pmp_7_addr_reg[19]_0 (\reg_pmp_7_addr_reg[19] ),
        .\reg_pmp_7_addr_reg[23]_0 (\reg_pmp_7_addr_reg[23] ),
        .\reg_pmp_7_addr_reg[28]_0 (\reg_pmp_7_addr_reg[28] ),
        .\reg_pmp_7_addr_reg[28]_1 (\reg_pmp_7_addr_reg[28]_0 ),
        .\reg_pmp_7_addr_reg[29]_0 (\reg_pmp_7_addr_reg[29] ),
        .\reg_pmp_7_addr_reg[29]_1 (\reg_pmp_7_addr_reg[29]_0 ),
        .\reg_pmp_7_addr_reg[29]_2 (\reg_pmp_7_addr_reg[29]_1 ),
        .\reg_pmp_7_addr_reg[29]_3 (\reg_pmp_7_addr_reg[29]_2 ),
        .\reg_pmp_7_cfg_a_reg[0]_0 (frontend_io_ptw_pmp_7_cfg_a[0]),
        .\reg_pmp_7_cfg_a_reg[0]_1 (\reg_pmp_7_cfg_a_reg[0] ),
        .\reg_pmp_7_cfg_a_reg[1]_0 (frontend_io_ptw_pmp_7_cfg_a[1]),
        .\reg_sbadaddr_reg[0]_0 (\reg_sbadaddr_reg[0] ),
        .\reg_sbadaddr_reg[30]_0 (\reg_sbadaddr_reg[30]_3 ),
        .\reg_sbadaddr_reg[39]_0 (\reg_sbadaddr_reg[39] ),
        .\reg_sbadaddr_reg[39]_1 (\reg_sbadaddr_reg[39]_0 ),
        .\reg_sbadaddr_reg[39]_2 (\reg_sbadaddr_reg[39]_1 ),
        .\reg_sbadaddr_reg[39]_3 (\reg_sbadaddr_reg[39]_2 ),
        .\reg_scause_reg[0]_0 (\reg_scause_reg[0] ),
        .\reg_scause_reg[0]_1 (\reg_scause_reg[0]_0 ),
        .\reg_scause_reg[1]_0 (\reg_scause_reg[1] ),
        .\reg_scause_reg[1]_1 (\reg_scause_reg[1]_0 ),
        .\reg_sepc_reg[12]_0 (\reg_sepc_reg[12] ),
        .\reg_sepc_reg[26]_0 (\reg_sepc_reg[26] ),
        .\reg_sptbr_mode_reg[3]_0 (frontend_io_ptw_ptbr_mode),
        .\reg_sptbr_ppn_reg[0]_0 (\reg_sptbr_ppn_reg[0] ),
        .\reg_sscratch_reg[0]_0 (\reg_sscratch_reg[0] ),
        .\reg_sscratch_reg[45]_0 ({\reg_sscratch_reg[45] [4],csr_io_bp_0_address,\reg_sscratch_reg[45] [3:0]}),
        .\reg_sscratch_reg[45]_1 (\reg_sscratch_reg[45]_0 ),
        .reg_wfi_reg_0(reg_wfi_reg),
        .resp_valid_0_reg(resp_valid_0_reg),
        .resp_valid_1_reg(resp_valid_1_reg),
        .\s1_pc_reg[1] (\s1_pc_reg[1] ),
        .\s1_pc_reg[26] (\s1_pc_reg[26] ),
        .\s1_pc_reg[31] (\s1_pc_reg[31] ),
        .\s1_pc_reg[39] (\s1_pc_reg[39]_0 ),
        .\s1_pc_reg[39]_0 (\s1_pc_reg[39]_6 ),
        .\s1_pc_reg[4] (\s1_pc_reg[4]_0 ),
        .\s1_pc_reg[4]_0 (\s1_pc_reg[4] ),
        .\s1_pc_reg[5] (\s1_pc_reg[5] ),
        .\s1_req_addr_reg[2] (\s1_req_addr_reg[2] ),
        .\s1_req_addr_reg[2]_0 (\s1_req_addr_reg[2]_0 ),
        .\s1_req_addr_reg[2]_1 (\s1_req_addr_reg[2]_1 ),
        .\s1_req_addr_reg[2]_2 (\s1_req_addr_reg[2]_2 ),
        .\s1_req_addr_reg[31] (\s1_req_addr_reg[31] ),
        .s1_req_phys_reg(s1_req_phys_reg),
        .s1_req_phys_reg_0(s1_req_phys_reg_0),
        .\s1_req_typ_reg[0] (\s1_req_typ_reg[0] ),
        .\s1_req_typ_reg[0]_0 (\s1_req_typ_reg[0]_0 ),
        .\s1_req_typ_reg[0]_1 (\s1_req_typ_reg[0]_1 ),
        .\s1_req_typ_reg[0]_2 (\s1_req_typ_reg[0]_2 ),
        .\s1_req_typ_reg[0]_3 (\s1_req_typ_reg[0]_3 ),
        .\s1_req_typ_reg[1] (\s1_req_typ_reg[1] ),
        .\s2_pc_reg[1] (\s2_pc_reg[1] ),
        .s2_replay(s2_replay),
        .\s2_req_addr_reg[31] (\s2_req_addr_reg[31] ),
        .s2_tlb_resp_cacheable_reg(s2_tlb_resp_cacheable_reg),
        .s2_valid_reg(s2_valid_reg),
        .\state_reg[0] (\state_reg[0]_2 ),
        .sys_reset_reg(sys_reset_reg),
        .sys_reset_reg_0(sys_reset_reg_1),
        .sys_reset_reg_1(sys_reset_reg_2),
        .target_reset(target_reset),
        .tile_auto_int_sync_xing_sinklzy_in_0_sync_0(tile_auto_int_sync_xing_sinklzy_in_0_sync_0),
        .tile_auto_int_sync_xing_sinklzy_in_0_sync_1(tile_auto_int_sync_xing_sinklzy_in_0_sync_1),
        .tile_auto_int_sync_xing_sinklzy_in_1_sync_0(tile_auto_int_sync_xing_sinklzy_in_1_sync_0),
        .tile_auto_int_sync_xing_sinklzy_in_2_sync_0(tile_auto_int_sync_xing_sinklzy_in_2_sync_0),
        .tlb_io_req_bits_sfence_bits_rs2(tlb_io_req_bits_sfence_bits_rs2),
        .\valid_reg[0] (\valid_reg[0] ),
        .\valid_reg[0]_0 (\valid_reg[0]_0 ),
        .\valid_reg[1] (\valid_reg[1] ),
        .\valid_reg[1]_0 (\valid_reg[1]_0 ),
        .\valid_reg[2] (\valid_reg[2] ),
        .\valid_reg[3] (\valid_reg[3]_2 ),
        .\valid_reg[3]_0 (\valid_reg[3]_3 ),
        .\valid_reg[3]_1 (\valid_reg[3]_4 ),
        .\valid_reg[4] (\valid_reg[4] ),
        .\wb_ctrl_csr_reg[0] (\wb_ctrl_csr_reg[0]_0 ),
        .\wb_ctrl_csr_reg[0]_0 (\wb_ctrl_csr_reg[0]_1 ),
        .\wb_ctrl_csr_reg[0]_1 (\wb_ctrl_csr_reg[0]_2 ),
        .\wb_ctrl_csr_reg[0]_2 (\wb_ctrl_csr_reg[0]_3 ),
        .\wb_ctrl_csr_reg[0]_3 (\wb_ctrl_csr_reg[0]_4 ),
        .\wb_ctrl_csr_reg[0]_4 (\wb_ctrl_csr_reg[0]_5 ),
        .\wb_ctrl_csr_reg[0]_5 (\wb_ctrl_csr_reg[0]_6 ),
        .\wb_ctrl_csr_reg[0]_6 (\wb_ctrl_csr_reg[0]_7 ),
        .\wb_ctrl_csr_reg[0]_7 (\wb_ctrl_csr_reg[0]_8 ),
        .\wb_ctrl_csr_reg[0]_8 (\wb_ctrl_csr_reg[0]_9 ),
        .\wb_ctrl_csr_reg[0]_9 (\wb_ctrl_csr_reg[0]_10 ),
        .\wb_ctrl_csr_reg[2] (\reg_sscratch_reg[59] ),
        .\wb_ctrl_csr_reg[2]_0 (\wb_ctrl_csr_reg[2]_0 ),
        .\wb_ctrl_csr_reg[2]_1 (_T_1396_reg_r1_0_31_0_5_i_44_n_0),
        .wb_ctrl_mem_reg(wb_ctrl_mem),
        .wb_ctrl_mem_reg_0(wb_ctrl_mem_reg_0),
        .\wb_ctrl_mem_type_reg[0] (\valid_reg[3]_1 ),
        .\wb_reg_cause_reg[0] (csr_io_bp_0_control_action),
        .\wb_reg_cause_reg[0]_0 (\wb_reg_cause_reg[0]_0 ),
        .\wb_reg_cause_reg[0]_1 (\wb_reg_cause_reg[0]_1 ),
        .\wb_reg_cause_reg[0]_10 (\wb_reg_cause_reg[0]_10 ),
        .\wb_reg_cause_reg[0]_11 (\wb_reg_cause_reg[0]_11 ),
        .\wb_reg_cause_reg[0]_12 (\wb_reg_cause_reg[0]_12 ),
        .\wb_reg_cause_reg[0]_13 (\wb_reg_cause_reg[0]_13 ),
        .\wb_reg_cause_reg[0]_14 (\wb_reg_cause_reg[0]_14 ),
        .\wb_reg_cause_reg[0]_2 (\wb_reg_cause_reg[0]_2 ),
        .\wb_reg_cause_reg[0]_3 (\wb_reg_cause_reg[0]_3 ),
        .\wb_reg_cause_reg[0]_4 (\wb_reg_cause_reg[0]_4 ),
        .\wb_reg_cause_reg[0]_5 (\wb_reg_cause_reg[0]_5 ),
        .\wb_reg_cause_reg[0]_6 (\wb_reg_cause_reg[0]_6 ),
        .\wb_reg_cause_reg[0]_7 (\wb_reg_cause_reg[0]_7 ),
        .\wb_reg_cause_reg[0]_8 (\wb_reg_cause_reg[0]_8 ),
        .\wb_reg_cause_reg[0]_9 (\wb_reg_cause_reg[0]_9 ),
        .\wb_reg_cause_reg[1] ({csr_n_747,csr_n_748}),
        .\wb_reg_cause_reg[2] (\wb_reg_cause_reg[2]_0 ),
        .\wb_reg_cause_reg[63] (\wb_reg_cause_reg[63]_0 ),
        .\wb_reg_cause_reg[63]_0 ({wb_reg_cause[63],wb_reg_cause[1:0]}),
        .\wb_reg_cause_reg[63]_1 (\wb_reg_cause_reg[63]_1 ),
        .\wb_reg_cause_reg[63]_2 (\wb_reg_cause_reg[63]_2 ),
        .\wb_reg_cause_reg[63]_3 (\wb_reg_cause_reg[63]_3 ),
        .\wb_reg_cause_reg[63]_4 (\wb_reg_cause_reg[63]_4 ),
        .\wb_reg_cause_reg[63]_5 (\wb_reg_cause_reg[63]_5 ),
        .\wb_reg_cause_reg[63]_6 (\wb_reg_cause_reg[63]_6 ),
        .wb_reg_flush_pipe(wb_reg_flush_pipe),
        .wb_reg_flush_pipe0(wb_reg_flush_pipe0),
        .\wb_reg_inst_reg[21] (\wb_reg_inst_reg[21]_0 ),
        .\wb_reg_inst_reg[21]_0 (\wb_reg_inst_reg[21]_1 ),
        .\wb_reg_inst_reg[21]_1 (\wb_reg_inst_reg[21]_2 ),
        .\wb_reg_inst_reg[21]_2 (\wb_reg_inst_reg[21]_3 ),
        .\wb_reg_inst_reg[21]_3 (\wb_reg_inst_reg[21]_4 ),
        .\wb_reg_inst_reg[21]_4 (\wb_reg_inst_reg[21]_5 ),
        .\wb_reg_inst_reg[21]_5 (\reg_scause_reg[3] ),
        .\wb_reg_inst_reg[22] (\wb_reg_inst_reg[22]_0 ),
        .\wb_reg_inst_reg[22]_0 (\reg_sptbr_ppn[19]_i_4_n_0 ),
        .\wb_reg_inst_reg[22]_1 (\wb_reg_inst_reg[22]_1 ),
        .\wb_reg_inst_reg[22]_2 (wb_reg_xcpt_i_2_n_0),
        .\wb_reg_inst_reg[26] (\wb_reg_inst_reg[26]_0 ),
        .\wb_reg_inst_reg[29] (\wb_reg_inst_reg[29]_0 ),
        .\wb_reg_inst_reg[29]_0 (\wb_reg_inst_reg[29]_1 ),
        .\wb_reg_inst_reg[30] (\wb_reg_inst_reg[30]_0 ),
        .\wb_reg_inst_reg[30]_0 (\wb_reg_inst_reg[30]_1 ),
        .\wb_reg_inst_reg[31] ({\reg_bp_0_control_tmatch_reg[1] [13:11],csr_io_rw_addr[8],\reg_bp_0_control_tmatch_reg[1] [10:9],csr_io_rw_addr[5],\reg_bp_0_control_tmatch_reg[1] [8],csr_io_rw_addr[3],\reg_bp_0_control_tmatch_reg[1] [7:5]}),
        .\wb_reg_pc_reg[39] ({\reg_dpc_reg[39] [38],\reg_dpc_reg[39] [0]}),
        .\wb_reg_pc_reg[39]_0 (\wb_reg_pc_reg[39]_1 ),
        .\wb_reg_pc_reg[39]_1 (\wb_reg_pc_reg[39]_2 ),
        .\wb_reg_pc_reg[39]_2 (\wb_reg_pc_reg[39]_3 ),
        .wb_reg_replay_reg(wb_reg_replay_reg_0),
        .wb_reg_replay_reg_0(wb_reg_replay_reg_1),
        .wb_reg_replay_reg_1(wb_reg_replay),
        .wb_reg_replay_reg_2(frontend_io_cpu_req_bits_speculative),
        .wb_reg_valid_reg(\valid_reg[3] ),
        .wb_reg_valid_reg_0(frontend_io_cpu_sfence_valid),
        .wb_reg_valid_reg_1(wb_reg_valid),
        .wb_reg_valid_reg_2(reg_debug_reg),
        .wb_reg_valid_reg_3(core__116_i_10_n_0),
        .wb_reg_valid_reg_4(\s1_pc[3]_i_7_n_0 ),
        .wb_reg_valid_reg_5(wb_reg_valid_reg_0),
        .wb_reg_xcpt0(wb_reg_xcpt0),
        .wb_reg_xcpt_reg(core__506_i_2_n_0),
        .wb_reg_xcpt_reg_0(wb_reg_xcpt));
  LUT4 #(
    .INIT(16'h00AE)) 
    data_arrays_0_0_reg_i_30
       (.I0(dcacheArb_io_requestor_1_req_valid),
        .I1(\state_reg[0]_0 ),
        .I2(\state_reg[1]_1 ),
        .I3(data_arrays_0_0_reg_i_53_n_0),
        .O(_T_481));
  LUT6 #(
    .INIT(64'h0C0D0C0D0C0B0C0C)) 
    data_arrays_0_0_reg_i_53
       (.I0(\s1_req_cmd_reg[4] [2]),
        .I1(\s1_req_cmd_reg[4] [4]),
        .I2(\state_reg[0]_1 ),
        .I3(\s1_req_cmd_reg[4] [3]),
        .I4(\s1_req_cmd_reg[4] [0]),
        .I5(\s1_req_cmd_reg[4] [1]),
        .O(data_arrays_0_0_reg_i_53_n_0));
  (* SOFT_HLUTNM = "soft_lutpair1863" *) 
  LUT4 #(
    .INIT(16'h00F8)) 
    dcache_blocked_i_1
       (.I0(ex_ctrl_mem),
        .I1(ex_reg_valid),
        .I2(dcache_blocked),
        .I3(dcacheArb_io_requestor_1_req_ready),
        .O(dcache_blocked0));
  FDRE #(
    .INIT(1'b0)) 
    dcache_blocked_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(dcache_blocked0),
        .Q(dcache_blocked),
        .R(\<const0> ));
  MulDiv div
       (.CO(CO),
        .D(\divisor_reg[57] [2:0]),
        .DI(DI),
        .O(O),
        .Q(ex_ctrl_alu_fn),
        .S(S),
        ._GEN_274(_GEN_274),
        ._T_1396__T_2475_addr({_T_1396__T_2475_addr,\ex_reg_rs_msb_1_reg[61]_1 }),
        ._T_1406(_T_1406_1),
        ._T_1416(_T_1416_0),
        ._T_2177(_T_2177),
        ._T_2222(_T_2222),
        ._T_2373(_T_2373),
        ._T_2518(_T_2518),
        .\_T_2547_reg[1] (\_T_2547_reg[1]_0 ),
        .\_T_2547_reg[31] (\_T_2547_reg[31]_0 ),
        .\_T_2547_reg[31]_0 (_T_2547[31:8]),
        .\_T_2547_reg[31]_1 ({_T_2549[31:17],\_T_2547_reg[16]_0 ,_T_2549[15:8]}),
        ._T_2770({_T_2770[20],_T_2770[17],_T_2770[14],_T_2770[9],_T_2770[6],_T_2770[1]}),
        .\buf__data_reg[14] (ibuf_n_64),
        .\buf__data_reg[2] (\buf__data_reg[2] ),
        .\buf__data_reg[3] (\buf__data_reg[3] ),
        .\buf__data_reg[4] (\buf__data_reg[4] ),
        .\bypass_mux_1_reg[32] ({\bypass_mux_1_reg_n_0_[32] ,\bypass_mux_1_reg_n_0_[31] ,\bypass_mux_1_reg_n_0_[30] ,\bypass_mux_1_reg_n_0_[29] ,\bypass_mux_1_reg_n_0_[28] ,\bypass_mux_1_reg_n_0_[27] ,\bypass_mux_1_reg_n_0_[26] ,\bypass_mux_1_reg_n_0_[25] ,\bypass_mux_1_reg_n_0_[24] ,\bypass_mux_1_reg_n_0_[23] ,\bypass_mux_1_reg_n_0_[22] ,\bypass_mux_1_reg_n_0_[21] ,\bypass_mux_1_reg_n_0_[20] ,\bypass_mux_1_reg_n_0_[19] ,\bypass_mux_1_reg_n_0_[18] ,\bypass_mux_1_reg_n_0_[17] ,\bypass_mux_1_reg_n_0_[16] ,\bypass_mux_1_reg_n_0_[15] ,\bypass_mux_1_reg_n_0_[14] ,\bypass_mux_1_reg_n_0_[13] ,\bypass_mux_1_reg_n_0_[12] ,\bypass_mux_1_reg_n_0_[11] ,\bypass_mux_1_reg_n_0_[10] ,\bypass_mux_1_reg_n_0_[9] ,\bypass_mux_1_reg_n_0_[8] ,\bypass_mux_1_reg_n_0_[7] ,\bypass_mux_1_reg_n_0_[6] ,\bypass_mux_1_reg_n_0_[5] ,\bypass_mux_1_reg_n_0_[4] ,\mem_reg_rs2_reg[3]_1 [1],\bypass_mux_1_reg_n_0_[2] ,\mem_reg_rs2_reg[3]_1 [0],\bypass_mux_1_reg_n_0_[0] }),
        .\bypass_mux_1_reg[33] (\bypass_mux_1_reg_n_0_[33] ),
        .\bypass_mux_1_reg[34] (\bypass_mux_1_reg_n_0_[34] ),
        .\bypass_mux_1_reg[35] (\bypass_mux_1_reg_n_0_[35] ),
        .\bypass_mux_1_reg[36] (\bypass_mux_1_reg_n_0_[36] ),
        .\bypass_mux_1_reg[37] (\bypass_mux_1_reg_n_0_[37] ),
        .\bypass_mux_1_reg[38] (\bypass_mux_2_reg[38]_0 ),
        .\bypass_mux_2_reg[0] (csr_n_664),
        .\bypass_mux_2_reg[0]_0 (\mem_reg_rs2_reg[0]_0 ),
        .\bypass_mux_2_reg[10] (\reg_mtvec_reg[10] ),
        .\bypass_mux_2_reg[11] (\reg_mtvec_reg[11] ),
        .\bypass_mux_2_reg[12] (\reg_mtvec_reg[12] ),
        .\bypass_mux_2_reg[13] (\reg_mtvec_reg[13] ),
        .\bypass_mux_2_reg[14] (\reg_mtvec_reg[14] ),
        .\bypass_mux_2_reg[15] (\reg_mtvec_reg[15] ),
        .\bypass_mux_2_reg[16] (\reg_mtvec_reg[16] ),
        .\bypass_mux_2_reg[17] (\reg_mtvec_reg[17] ),
        .\bypass_mux_2_reg[18] (\reg_mtvec_reg[18] ),
        .\bypass_mux_2_reg[19] (\reg_mtvec_reg[19] ),
        .\bypass_mux_2_reg[1] (csr_n_665),
        .\bypass_mux_2_reg[1]_0 (\mem_reg_rs2_reg[1]_0 ),
        .\bypass_mux_2_reg[20] (\reg_mtvec_reg[20]_0 ),
        .\bypass_mux_2_reg[21] (\reg_mtvec_reg[21]_0 ),
        .\bypass_mux_2_reg[22] (\reg_mtvec_reg[22]_0 ),
        .\bypass_mux_2_reg[23] (\reg_mtvec_reg[23] ),
        .\bypass_mux_2_reg[24] (\reg_mtvec_reg[24] ),
        .\bypass_mux_2_reg[25] (\reg_mtvec_reg[25] ),
        .\bypass_mux_2_reg[26] (\reg_mtvec_reg[26] ),
        .\bypass_mux_2_reg[27] (\reg_mtvec_reg[27] ),
        .\bypass_mux_2_reg[28] (\reg_mtvec_reg[28] ),
        .\bypass_mux_2_reg[29] (\reg_mtvec_reg[29]_7 ),
        .\bypass_mux_2_reg[2] (csr_n_666),
        .\bypass_mux_2_reg[2]_0 (\mem_reg_rs2_reg[2]_0 ),
        .\bypass_mux_2_reg[30] (csr_n_678),
        .\bypass_mux_2_reg[30]_0 (\reg_mtvec_reg[30] ),
        .\bypass_mux_2_reg[31] (csr_n_677),
        .\bypass_mux_2_reg[31]_0 (\reg_mtvec_reg[31] ),
        .\bypass_mux_2_reg[32] (csr_n_676),
        .\bypass_mux_2_reg[32]_0 (\reg_stvec_reg[32] ),
        .\bypass_mux_2_reg[33] (csr_n_675),
        .\bypass_mux_2_reg[33]_0 (\reg_stvec_reg[33] ),
        .\bypass_mux_2_reg[34] (csr_n_674),
        .\bypass_mux_2_reg[34]_0 (\reg_stvec_reg[34] ),
        .\bypass_mux_2_reg[35] (csr_n_673),
        .\bypass_mux_2_reg[35]_0 (\reg_stvec_reg[35] ),
        .\bypass_mux_2_reg[36] (csr_n_672),
        .\bypass_mux_2_reg[36]_0 (\reg_stvec_reg[36] ),
        .\bypass_mux_2_reg[37] (csr_n_671),
        .\bypass_mux_2_reg[37]_0 (\reg_stvec_reg[37] ),
        .\bypass_mux_2_reg[38] (csr_n_670),
        .\bypass_mux_2_reg[38]_0 (\reg_stvec_reg[38] ),
        .\bypass_mux_2_reg[39] (csr_n_702),
        .\bypass_mux_2_reg[39]_0 (\reg_sscratch_reg[62] [0]),
        .\bypass_mux_2_reg[3] (csr_n_667),
        .\bypass_mux_2_reg[3]_0 (\mem_reg_rs2_reg[3]_0 ),
        .\bypass_mux_2_reg[40] (csr_n_701),
        .\bypass_mux_2_reg[40]_0 (\reg_sscratch_reg[62] [1]),
        .\bypass_mux_2_reg[41] (csr_n_700),
        .\bypass_mux_2_reg[41]_0 (\reg_sscratch_reg[62] [2]),
        .\bypass_mux_2_reg[42] (csr_n_699),
        .\bypass_mux_2_reg[42]_0 (\reg_sscratch_reg[62] [3]),
        .\bypass_mux_2_reg[43] (csr_n_698),
        .\bypass_mux_2_reg[43]_0 (\reg_sscratch_reg[62] [4]),
        .\bypass_mux_2_reg[44] (csr_n_689),
        .\bypass_mux_2_reg[44]_0 (\reg_sscratch_reg[62] [5]),
        .\bypass_mux_2_reg[45] (csr_n_697),
        .\bypass_mux_2_reg[45]_0 (\reg_sscratch_reg[62] [6]),
        .\bypass_mux_2_reg[46] (csr_n_696),
        .\bypass_mux_2_reg[46]_0 (\reg_sscratch_reg[62] [7]),
        .\bypass_mux_2_reg[47] (csr_n_688),
        .\bypass_mux_2_reg[47]_0 (\reg_sscratch_reg[62] [8]),
        .\bypass_mux_2_reg[48] (csr_n_687),
        .\bypass_mux_2_reg[48]_0 (\reg_sscratch_reg[62] [9]),
        .\bypass_mux_2_reg[49] (csr_n_686),
        .\bypass_mux_2_reg[49]_0 (\reg_sscratch_reg[62] [10]),
        .\bypass_mux_2_reg[4] (csr_n_668),
        .\bypass_mux_2_reg[4]_0 (\mem_reg_rs2_reg[4]_0 ),
        .\bypass_mux_2_reg[50] (csr_n_685),
        .\bypass_mux_2_reg[50]_0 (\reg_sscratch_reg[62] [11]),
        .\bypass_mux_2_reg[51] (csr_n_684),
        .\bypass_mux_2_reg[51]_0 (\reg_sscratch_reg[62] [12]),
        .\bypass_mux_2_reg[52] (csr_n_683),
        .\bypass_mux_2_reg[52]_0 (\reg_sscratch_reg[62] [13]),
        .\bypass_mux_2_reg[53] (csr_n_695),
        .\bypass_mux_2_reg[53]_0 (\reg_sscratch_reg[62] [14]),
        .\bypass_mux_2_reg[54] (csr_n_694),
        .\bypass_mux_2_reg[54]_0 (\reg_sscratch_reg[62] [15]),
        .\bypass_mux_2_reg[55] (csr_n_693),
        .\bypass_mux_2_reg[55]_0 (\reg_sscratch_reg[62] [16]),
        .\bypass_mux_2_reg[56] (csr_n_682),
        .\bypass_mux_2_reg[56]_0 (\reg_sscratch_reg[62] [17]),
        .\bypass_mux_2_reg[57] (csr_n_681),
        .\bypass_mux_2_reg[57]_0 (\reg_sscratch_reg[62] [18]),
        .\bypass_mux_2_reg[58] (csr_n_680),
        .\bypass_mux_2_reg[58]_0 (\reg_sscratch_reg[62] [19]),
        .\bypass_mux_2_reg[59] (csr_n_703),
        .\bypass_mux_2_reg[59]_0 (\reg_sscratch_reg[62] [20]),
        .\bypass_mux_2_reg[5] (csr_n_669),
        .\bypass_mux_2_reg[5]_0 (\mem_reg_rs2_reg[5]_0 ),
        .\bypass_mux_2_reg[60] (csr_n_692),
        .\bypass_mux_2_reg[60]_0 (\reg_sscratch_reg[62] [21]),
        .\bypass_mux_2_reg[61] (csr_n_691),
        .\bypass_mux_2_reg[61]_0 (\reg_sscratch_reg[62] [22]),
        .\bypass_mux_2_reg[62] (csr_n_690),
        .\bypass_mux_2_reg[62]_0 (\reg_sscratch_reg[62] [23]),
        .\bypass_mux_2_reg[63] (csr_n_679),
        .\bypass_mux_2_reg[6] (csr_n_642),
        .\bypass_mux_2_reg[6]_0 (\mem_reg_rs2_reg[6]_0 ),
        .\bypass_mux_2_reg[7] (csr_n_641),
        .\bypass_mux_2_reg[7]_0 (\mem_reg_rs2_reg[7]_0 ),
        .\bypass_mux_2_reg[8] (csr_n_643),
        .\bypass_mux_2_reg[8]_0 (\reg_mtvec_reg[8] ),
        .\bypass_mux_2_reg[9] (csr_n_644),
        .\bypass_mux_2_reg[9]_0 (reg_mip_seip_reg_0),
        .\bypass_mux_2_reg[9]_1 (\bypass_mux_2_reg[9]_0 ),
        .\count_reg[0]_0 (\count_reg[0] ),
        .dcacheArb_io_requestor_1_ordered(dcacheArb_io_requestor_1_ordered),
        .dcacheArb_io_requestor_1_replay_next(dcacheArb_io_requestor_1_replay_next),
        .dcacheArb_io_requestor_1_req_ready(dcacheArb_io_requestor_1_req_ready),
        .dcacheArb_io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),
        .dcacheArb_io_requestor_1_resp_bits_data(dcacheArb_io_requestor_1_resp_bits_data),
        .dcacheArb_io_requestor_1_resp_bits_data_word_bypass(dcacheArb_io_requestor_1_resp_bits_data_word_bypass),
        .dcacheArb_io_requestor_1_resp_bits_replay(dcacheArb_io_requestor_1_resp_bits_replay),
        .dcacheArb_io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),
        .dcacheArb_io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),
        .\divisor_reg[10]_0 (div_n_219),
        .\divisor_reg[11]_0 (div_n_220),
        .\divisor_reg[12]_0 (div_n_221),
        .\divisor_reg[13]_0 (div_n_222),
        .\divisor_reg[14]_0 (div_n_223),
        .\divisor_reg[15]_0 (div_n_224),
        .\divisor_reg[15]_1 (\divisor_reg[15] ),
        .\divisor_reg[15]_10 (\divisor_reg[15]_8 ),
        .\divisor_reg[15]_2 (\divisor_reg[15]_0 ),
        .\divisor_reg[15]_3 (\divisor_reg[15]_1 ),
        .\divisor_reg[15]_4 (\divisor_reg[15]_2 ),
        .\divisor_reg[15]_5 (\divisor_reg[15]_3 ),
        .\divisor_reg[15]_6 (\divisor_reg[15]_4 ),
        .\divisor_reg[15]_7 (\divisor_reg[15]_5 ),
        .\divisor_reg[15]_8 (\divisor_reg[15]_6 ),
        .\divisor_reg[15]_9 (\divisor_reg[15]_7 ),
        .\divisor_reg[18]_0 (div_n_225),
        .\divisor_reg[18]_1 (\divisor_reg[18] ),
        .\divisor_reg[19]_0 (div_n_226),
        .\divisor_reg[1]_0 (\divisor_reg[1] ),
        .\divisor_reg[20]_0 (div_n_227),
        .\divisor_reg[21]_0 (div_n_228),
        .\divisor_reg[22]_0 (div_n_229),
        .\divisor_reg[23]_0 (div_n_230),
        .\divisor_reg[25]_0 (\divisor_reg[57] [3]),
        .\divisor_reg[32]_0 (\divisor_reg[32] ),
        .\divisor_reg[32]_1 (\divisor_reg[32]_0 ),
        .\divisor_reg[32]_2 (\divisor_reg[32]_1 ),
        .\divisor_reg[35]_0 (\divisor_reg[35] ),
        .\divisor_reg[50]_0 (div_n_234),
        .\divisor_reg[51]_0 (div_n_235),
        .\divisor_reg[51]_1 (\divisor_reg[51] ),
        .\divisor_reg[52]_0 (div_n_236),
        .\divisor_reg[52]_1 (\divisor_reg[52] ),
        .\divisor_reg[53]_0 (div_n_237),
        .\divisor_reg[54]_0 (div_n_238),
        .\divisor_reg[55]_0 (div_n_239),
        .\divisor_reg[57]_0 (\divisor_reg[57] [5:4]),
        .\divisor_reg[8]_0 (div_n_218),
        .doUncachedResp_reg(doUncachedResp_reg),
        .ex_ctrl_alu_dw_reg(req_dw_reg),
        .ex_ctrl_div_reg(ex_ctrl_div),
        .ex_ctrl_mem(ex_ctrl_mem),
        .ex_ctrl_mem_reg(div_n_368),
        .ex_ctrl_mem_reg_0(ex_ctrl_mem_reg_1),
        .\ex_reg_inst_reg[11] (\mem_reg_inst_reg[31]_0 [4:0]),
        .ex_reg_load_use(ex_reg_load_use),
        .ex_reg_replay(ex_reg_replay),
        .ex_reg_rs_bypass_0_reg(ex_reg_rs_bypass_0_reg_0),
        .ex_reg_rs_bypass_1(ex_reg_rs_bypass_1),
        .\ex_reg_rs_lsb_0_reg[1] (\ex_reg_rs_lsb_0_reg[1]_0 ),
        .\ex_reg_rs_lsb_0_reg[1]_0 (ex_reg_rs_lsb_0),
        .\ex_reg_rs_lsb_1_reg[1] ({\ex_reg_rs_lsb_1_reg_n_0_[1] ,\ex_reg_rs_lsb_1_reg_n_0_[0] }),
        .\ex_reg_rs_msb_0_reg[27] (\ex_reg_rs_msb_0_reg[27]_0 ),
        .\ex_reg_rs_msb_0_reg[61] ({\ex_reg_rs_msb_0_reg_n_0_[61] ,\ex_reg_rs_msb_0_reg_n_0_[60] ,\ex_reg_rs_msb_0_reg_n_0_[59] ,\ex_reg_rs_msb_0_reg_n_0_[58] ,\ex_reg_rs_msb_0_reg_n_0_[57] ,\ex_reg_rs_msb_0_reg_n_0_[56] ,\ex_reg_rs_msb_0_reg_n_0_[55] ,\ex_reg_rs_msb_0_reg_n_0_[54] ,\ex_reg_rs_msb_0_reg_n_0_[53] ,\ex_reg_rs_msb_0_reg_n_0_[52] ,\ex_reg_rs_msb_0_reg_n_0_[51] ,\ex_reg_rs_msb_0_reg_n_0_[50] ,\ex_reg_rs_msb_0_reg_n_0_[49] ,\ex_reg_rs_msb_0_reg_n_0_[48] ,\ex_reg_rs_msb_0_reg_n_0_[47] ,\ex_reg_rs_msb_0_reg_n_0_[46] ,\ex_reg_rs_msb_0_reg_n_0_[45] ,\ex_reg_rs_msb_0_reg_n_0_[44] ,\ex_reg_rs_msb_0_reg_n_0_[43] ,\ex_reg_rs_msb_0_reg_n_0_[42] ,\ex_reg_rs_msb_0_reg_n_0_[41] ,\ex_reg_rs_msb_0_reg_n_0_[40] ,\ex_reg_rs_msb_0_reg_n_0_[39] ,\ex_reg_rs_msb_0_reg_n_0_[38] ,\ex_reg_rs_msb_0_reg_n_0_[37] ,\ex_reg_rs_msb_0_reg_n_0_[36] ,\ex_reg_rs_msb_0_reg_n_0_[35] ,\ex_reg_rs_msb_0_reg_n_0_[34] ,\ex_reg_rs_msb_0_reg_n_0_[33] ,\ex_reg_rs_msb_0_reg_n_0_[32] ,\ex_reg_rs_msb_0_reg_n_0_[31] ,\ex_reg_rs_msb_0_reg_n_0_[30] ,\ex_reg_rs_msb_0_reg_n_0_[29] ,\ex_reg_rs_msb_0_reg_n_0_[28] ,\ex_reg_rs_msb_0_reg_n_0_[27] ,\ex_reg_rs_msb_0_reg_n_0_[26] ,\ex_reg_rs_msb_0_reg_n_0_[25] ,\ex_reg_rs_msb_0_reg_n_0_[24] ,\ex_reg_rs_msb_0_reg_n_0_[23] ,\ex_reg_rs_msb_0_reg_n_0_[22] ,\ex_reg_rs_msb_0_reg_n_0_[21] ,\ex_reg_rs_msb_0_reg_n_0_[20] ,\ex_reg_rs_msb_0_reg_n_0_[19] ,\ex_reg_rs_msb_0_reg_n_0_[18] ,\ex_reg_rs_msb_0_reg_n_0_[17] ,\ex_reg_rs_msb_0_reg_n_0_[16] ,\ex_reg_rs_msb_0_reg_n_0_[15] ,\ex_reg_rs_msb_0_reg_n_0_[14] ,\ex_reg_rs_msb_0_reg_n_0_[13] ,\ex_reg_rs_msb_0_reg_n_0_[12] ,\ex_reg_rs_msb_0_reg_n_0_[11] ,\ex_reg_rs_msb_0_reg_n_0_[10] ,\ex_reg_rs_msb_0_reg_n_0_[9] ,\ex_reg_rs_msb_0_reg_n_0_[8] ,\ex_reg_rs_msb_0_reg_n_0_[7] ,\ex_reg_rs_msb_0_reg_n_0_[6] ,\ex_reg_rs_msb_0_reg_n_0_[5] ,\ex_reg_rs_msb_0_reg_n_0_[4] ,\ex_reg_rs_msb_0_reg_n_0_[3] ,\ex_reg_rs_msb_0_reg_n_0_[2] ,\ex_reg_rs_msb_0_reg_n_0_[1] ,\ex_reg_rs_msb_0_reg_n_0_[0] }),
        .\ex_reg_rs_msb_1_reg[29] (\ex_reg_rs_msb_1_reg[29]_0 ),
        .\ex_reg_rs_msb_1_reg[61] (_T_1856),
        .\ex_reg_rs_msb_1_reg[61]_0 (\ex_reg_rs_msb_1_reg[61]_0 ),
        .\ex_reg_rs_msb_1_reg[61]_1 (\ex_reg_rs_msb_1_reg[61]_2 ),
        .\ex_reg_rs_msb_1_reg[61]_2 ({\ex_reg_rs_msb_1_reg_n_0_[61] ,\ex_reg_rs_msb_1_reg_n_0_[60] ,\ex_reg_rs_msb_1_reg_n_0_[59] ,\ex_reg_rs_msb_1_reg_n_0_[58] ,\ex_reg_rs_msb_1_reg_n_0_[57] ,\ex_reg_rs_msb_1_reg_n_0_[56] ,\ex_reg_rs_msb_1_reg_n_0_[55] ,\ex_reg_rs_msb_1_reg_n_0_[54] ,\ex_reg_rs_msb_1_reg_n_0_[53] ,\ex_reg_rs_msb_1_reg_n_0_[52] ,\ex_reg_rs_msb_1_reg_n_0_[51] ,\ex_reg_rs_msb_1_reg_n_0_[50] ,\ex_reg_rs_msb_1_reg_n_0_[49] ,\ex_reg_rs_msb_1_reg_n_0_[48] ,\ex_reg_rs_msb_1_reg_n_0_[47] ,\ex_reg_rs_msb_1_reg_n_0_[46] ,\ex_reg_rs_msb_1_reg_n_0_[45] ,\ex_reg_rs_msb_1_reg_n_0_[44] ,\ex_reg_rs_msb_1_reg_n_0_[43] ,\ex_reg_rs_msb_1_reg_n_0_[42] ,\ex_reg_rs_msb_1_reg_n_0_[41] ,\ex_reg_rs_msb_1_reg_n_0_[40] ,\ex_reg_rs_msb_1_reg_n_0_[39] ,\ex_reg_rs_msb_1_reg_n_0_[38] ,\ex_reg_rs_msb_1_reg_n_0_[37] ,\ex_reg_rs_msb_1_reg_n_0_[36] ,\ex_reg_rs_msb_1_reg_n_0_[35] ,\ex_reg_rs_msb_1_reg_n_0_[34] ,\ex_reg_rs_msb_1_reg_n_0_[33] ,\ex_reg_rs_msb_1_reg_n_0_[32] ,\ex_reg_rs_msb_1_reg_n_0_[31] ,\ex_reg_rs_msb_1_reg_n_0_[30] ,\ex_reg_rs_msb_1_reg_n_0_[29] ,\ex_reg_rs_msb_1_reg_n_0_[28] ,\ex_reg_rs_msb_1_reg_n_0_[27] ,\ex_reg_rs_msb_1_reg_n_0_[26] ,\ex_reg_rs_msb_1_reg_n_0_[25] ,\ex_reg_rs_msb_1_reg_n_0_[24] ,\ex_reg_rs_msb_1_reg_n_0_[23] ,\ex_reg_rs_msb_1_reg_n_0_[22] ,\ex_reg_rs_msb_1_reg_n_0_[21] ,\ex_reg_rs_msb_1_reg_n_0_[20] ,\ex_reg_rs_msb_1_reg_n_0_[19] ,\ex_reg_rs_msb_1_reg_n_0_[18] ,\ex_reg_rs_msb_1_reg_n_0_[17] ,\ex_reg_rs_msb_1_reg_n_0_[16] ,\ex_reg_rs_msb_1_reg_n_0_[15] ,\ex_reg_rs_msb_1_reg_n_0_[14] ,\ex_reg_rs_msb_1_reg_n_0_[13] ,\ex_reg_rs_msb_1_reg_n_0_[12] ,\ex_reg_rs_msb_1_reg_n_0_[11] ,\ex_reg_rs_msb_1_reg_n_0_[10] ,\ex_reg_rs_msb_1_reg_n_0_[9] ,\ex_reg_rs_msb_1_reg_n_0_[8] ,\ex_reg_rs_msb_1_reg_n_0_[7] ,\ex_reg_rs_msb_1_reg_n_0_[6] ,\ex_reg_rs_msb_1_reg_n_0_[5] ,\ex_reg_rs_msb_1_reg_n_0_[4] ,\ex_reg_rs_msb_1_reg_n_0_[3] ,\ex_reg_rs_msb_1_reg_n_0_[2] ,\ex_reg_rs_msb_1_reg_n_0_[1] ,\ex_reg_rs_msb_1_reg_n_0_[0] }),
        .ex_reg_valid_reg(ex_reg_valid),
        .host_clk(host_clk),
        .ibuf_io_inst_0_bits_inst_rs2({ibuf_io_inst_0_bits_inst_rs2[2],ibuf_io_inst_0_bits_inst_rs2[0]}),
        .id_reg_fence_reg(id_reg_fence_reg_0),
        .mem_ctrl_wxd(mem_ctrl_wxd),
        .mem_reg_replay0(mem_reg_replay0),
        .mem_reg_rs2({mem_reg_rs2[63:58],mem_reg_rs2[56],mem_reg_rs2[49:42],mem_reg_rs2[40:26],mem_reg_rs2[24],mem_reg_rs2[17:16],mem_reg_rs2[5:2],mem_reg_rs2[0]}),
        .\mem_reg_rs2_reg[25] (\mem_reg_rs2_reg[25]_0 ),
        .mem_reg_valid_reg(mem_reg_valid_reg_0),
        .mem_reg_valid_reg_0(mem_reg_replay_reg_0),
        .mem_reg_valid_reg_1(mem_reg_valid),
        .mem_reg_xcpt_reg(mem_reg_xcpt),
        .nBufValid_reg(nBufValid_reg_3),
        .nBufValid_reg_0(ibuf_n_56),
        .neg_out_reg_0(neg_out_reg),
        .neg_out_reg_1(div_n_526),
        .p_0_in32_out(p_31_in),
        .\remainder_reg[0]_0 (div_n_240),
        .\remainder_reg[103]_0 (\remainder_reg[103] ),
        .\remainder_reg[103]_1 (\remainder_reg[103]_0 ),
        .\remainder_reg[103]_2 (\remainder_reg[103]_1 ),
        .\remainder_reg[103]_3 (\remainder_reg[103]_2 ),
        .\remainder_reg[107]_0 (\remainder_reg[107] ),
        .\remainder_reg[107]_1 (\remainder_reg[107]_0 ),
        .\remainder_reg[107]_2 (\remainder_reg[107]_1 ),
        .\remainder_reg[10]_0 (div_n_147),
        .\remainder_reg[111]_0 (\remainder_reg[111] ),
        .\remainder_reg[111]_1 (\remainder_reg[111]_0 ),
        .\remainder_reg[111]_2 (\remainder_reg[111]_1 ),
        .\remainder_reg[115]_0 (\remainder_reg[115] ),
        .\remainder_reg[115]_1 (\remainder_reg[115]_0 ),
        .\remainder_reg[115]_2 (\remainder_reg[115]_1 ),
        .\remainder_reg[115]_3 (\remainder_reg[115]_2 ),
        .\remainder_reg[119]_0 (\remainder_reg[119] ),
        .\remainder_reg[119]_1 (\remainder_reg[119]_0 ),
        .\remainder_reg[11]_0 (div_n_148),
        .\remainder_reg[123]_0 (\remainder_reg[123] ),
        .\remainder_reg[123]_1 (\remainder_reg[123]_0 ),
        .\remainder_reg[127]_0 (\remainder_reg[127] ),
        .\remainder_reg[127]_1 (\remainder_reg[127]_0 ),
        .\remainder_reg[127]_2 (\remainder_reg[127]_1 ),
        .\remainder_reg[127]_3 (\remainder_reg[127]_2 ),
        .\remainder_reg[127]_4 (\remainder_reg[127]_3 ),
        .\remainder_reg[127]_5 (\remainder_reg[127]_4 ),
        .\remainder_reg[127]_6 (\remainder_reg[127]_5 ),
        .\remainder_reg[127]_7 (\remainder_reg[127]_6 ),
        .\remainder_reg[127]_8 (\remainder_reg[127]_7 ),
        .\remainder_reg[128]_0 (\remainder_reg[128] ),
        .\remainder_reg[129]_0 (\remainder_reg[129] ),
        .\remainder_reg[129]_1 (\remainder_reg[129]_0 ),
        .\remainder_reg[129]_2 (_T_216),
        .\remainder_reg[129]_3 (\remainder_reg[129]_1 ),
        .\remainder_reg[12]_0 (div_n_149),
        .\remainder_reg[13]_0 (div_n_150),
        .\remainder_reg[14]_0 (div_n_151),
        .\remainder_reg[15]_0 (div_n_152),
        .\remainder_reg[16]_0 (div_n_153),
        .\remainder_reg[17]_0 (div_n_154),
        .\remainder_reg[18]_0 (div_n_155),
        .\remainder_reg[19]_0 (div_n_156),
        .\remainder_reg[1]_0 (div_n_138),
        .\remainder_reg[20]_0 (div_n_157),
        .\remainder_reg[21]_0 (div_n_158),
        .\remainder_reg[22]_0 (div_n_159),
        .\remainder_reg[23]_0 (div_n_160),
        .\remainder_reg[24]_0 (div_n_161),
        .\remainder_reg[25]_0 (div_n_162),
        .\remainder_reg[26]_0 (div_n_163),
        .\remainder_reg[27]_0 (div_n_164),
        .\remainder_reg[28]_0 (div_n_165),
        .\remainder_reg[29]_0 (div_n_166),
        .\remainder_reg[2]_0 (div_n_139),
        .\remainder_reg[30]_0 (div_n_167),
        .\remainder_reg[31]_0 (\remainder_reg[31] ),
        .\remainder_reg[32]_0 (div_n_170),
        .\remainder_reg[33]_0 (\remainder_reg[33] ),
        .\remainder_reg[33]_1 (\remainder_reg[33]_0 ),
        .\remainder_reg[34]_0 (\remainder_reg[34] ),
        .\remainder_reg[34]_1 (\remainder_reg[34]_0 ),
        .\remainder_reg[35]_0 (\remainder_reg[35] ),
        .\remainder_reg[35]_1 (\remainder_reg[35]_0 ),
        .\remainder_reg[36]_0 (\remainder_reg[36] ),
        .\remainder_reg[36]_1 (\remainder_reg[36]_0 ),
        .\remainder_reg[37]_0 (\remainder_reg[37] ),
        .\remainder_reg[37]_1 (\remainder_reg[37]_0 ),
        .\remainder_reg[38]_0 (\remainder_reg[38] ),
        .\remainder_reg[38]_1 (\remainder_reg[38]_0 ),
        .\remainder_reg[39]_0 (\remainder_reg[39] ),
        .\remainder_reg[39]_1 (\s1_req_addr_reg[39] [0]),
        .\remainder_reg[3]_0 (div_n_140),
        .\remainder_reg[41]_0 (\remainder_reg[41] ),
        .\remainder_reg[41]_1 (\s1_req_addr_reg[39] [1]),
        .\remainder_reg[42]_0 (\remainder_reg[42] ),
        .\remainder_reg[42]_1 (\s1_req_addr_reg[39] [2]),
        .\remainder_reg[43]_0 (\remainder_reg[43] ),
        .\remainder_reg[43]_1 (\s1_req_addr_reg[39] [3]),
        .\remainder_reg[44]_0 (\remainder_reg[44] ),
        .\remainder_reg[44]_1 (\s1_req_addr_reg[39] [4]),
        .\remainder_reg[46]_0 (\remainder_reg[46] ),
        .\remainder_reg[46]_1 (\s1_req_addr_reg[39] [5]),
        .\remainder_reg[47]_0 (\remainder_reg[47] ),
        .\remainder_reg[47]_1 (\s1_req_addr_reg[39] [6]),
        .\remainder_reg[49]_0 (\remainder_reg[49] ),
        .\remainder_reg[49]_1 (\s1_req_addr_reg[39] [7]),
        .\remainder_reg[4]_0 (div_n_141),
        .\remainder_reg[50]_0 (\remainder_reg[50] ),
        .\remainder_reg[50]_1 (\s1_req_addr_reg[39] [8]),
        .\remainder_reg[51]_0 (\remainder_reg[51] ),
        .\remainder_reg[51]_1 (\s1_req_addr_reg[39] [9]),
        .\remainder_reg[52]_0 (\remainder_reg[52] ),
        .\remainder_reg[52]_1 (\s1_req_addr_reg[39] [10]),
        .\remainder_reg[54]_0 (\remainder_reg[54] ),
        .\remainder_reg[54]_1 (\s1_req_addr_reg[39] [11]),
        .\remainder_reg[55]_0 (\remainder_reg[55] ),
        .\remainder_reg[55]_1 (\s1_req_addr_reg[39] [12]),
        .\remainder_reg[57]_0 (\remainder_reg[57] ),
        .\remainder_reg[57]_1 (\s1_req_addr_reg[39] [13]),
        .\remainder_reg[58]_0 (\remainder_reg[58] ),
        .\remainder_reg[58]_1 (\s1_req_addr_reg[39] [14]),
        .\remainder_reg[59]_0 (\remainder_reg[59] ),
        .\remainder_reg[5]_0 (div_n_142),
        .\remainder_reg[60]_0 (\remainder_reg[60] ),
        .\remainder_reg[60]_1 (\s1_req_addr_reg[39] [15]),
        .\remainder_reg[61]_0 (\remainder_reg[61] ),
        .\remainder_reg[61]_1 (\s1_req_addr_reg[39] [16]),
        .\remainder_reg[62]_0 (\remainder_reg[62] ),
        .\remainder_reg[62]_1 (\s1_req_addr_reg[39] [17]),
        .\remainder_reg[62]_2 (\remainder_reg[62]_0 ),
        .\remainder_reg[63]_0 (\remainder_reg[63] ),
        .\remainder_reg[64]_0 (\remainder_reg[64] ),
        .\remainder_reg[64]_1 (\remainder_reg[64]_0 ),
        .\remainder_reg[64]_10 (\remainder_reg[64]_9 ),
        .\remainder_reg[64]_2 (\remainder_reg[64]_1 ),
        .\remainder_reg[64]_3 (\remainder_reg[64]_2 ),
        .\remainder_reg[64]_4 (\remainder_reg[64]_3 ),
        .\remainder_reg[64]_5 (\remainder_reg[64]_4 ),
        .\remainder_reg[64]_6 (\remainder_reg[64]_5 ),
        .\remainder_reg[64]_7 (\remainder_reg[64]_6 ),
        .\remainder_reg[64]_8 (\remainder_reg[64]_7 ),
        .\remainder_reg[64]_9 (\remainder_reg[64]_8 ),
        .\remainder_reg[65]_0 (\remainder_reg[65] ),
        .\remainder_reg[6]_0 (div_n_143),
        .\remainder_reg[71]_0 (\remainder_reg[71] ),
        .\remainder_reg[75]_0 (\remainder_reg[75] ),
        .\remainder_reg[79]_0 (\remainder_reg[79] ),
        .\remainder_reg[7]_0 (div_n_144),
        .\remainder_reg[83]_0 (\remainder_reg[83] ),
        .\remainder_reg[87]_0 (\remainder_reg[87] ),
        .\remainder_reg[8]_0 (div_n_145),
        .\remainder_reg[91]_0 (\remainder_reg[91] ),
        .\remainder_reg[91]_1 (\remainder_reg[91]_0 ),
        .\remainder_reg[95]_0 (\remainder_reg[95] ),
        .\remainder_reg[95]_1 (\remainder_reg[95]_0 ),
        .\remainder_reg[99]_0 (\remainder_reg[99] ),
        .\remainder_reg[99]_1 (\remainder_reg[99]_0 ),
        .\remainder_reg[9]_0 (div_n_146),
        .\req_tag_reg[0]_0 (\req_tag_reg[0] ),
        .\req_tag_reg[0]_1 (\req_tag_reg[0]_0 ),
        .\req_tag_reg[1]_0 (\req_tag_reg[1]_4 ),
        .\req_tag_reg[1]_1 (\req_tag_reg[1] ),
        .\req_tag_reg[1]_2 (\req_tag_reg[1]_0 ),
        .\req_tag_reg[1]_3 (\req_tag_reg[1]_1 ),
        .\req_tag_reg[1]_4 (\req_tag_reg[1]_2 ),
        .\req_tag_reg[1]_5 (\req_tag_reg[1]_3 ),
        .\req_tag_reg[4]_0 (\req_tag_reg[4] ),
        .resHi_reg_0(resHi_reg),
        .\s2_req_cmd_reg[1] (\s2_req_cmd_reg[1] ),
        .\s2_req_tag_reg[5] (\s2_req_tag_reg[5]_0 ),
        .\s2_req_tag_reg[6] (\s2_req_tag_reg[6] ),
        .\s2_req_typ_reg[0] (\s2_req_typ_reg[0] ),
        .\state_reg[0]_0 (\state_reg[0] ),
        .\state_reg[1]_0 (\state_reg[1]_0 ),
        .\state_reg[2]_0 (\state_reg[2] ),
        .sys_reset_reg(sys_reset_reg_0),
        .target_reset(target_reset),
        .wb_ctrl_mem_reg(wb_ctrl_mem),
        .wb_ctrl_wxd_reg(wb_ctrl_wxd),
        .wb_reg_flush_pipe(wb_reg_flush_pipe),
        .\wb_reg_inst_reg[10] (\_T_2547[23]_i_3_n_0 ),
        .\wb_reg_inst_reg[11] (\reg_bp_0_control_tmatch_reg[1] [4:0]),
        .\wb_reg_inst_reg[11]_0 (\_T_2547[15]_i_3_n_0 ),
        .\wb_reg_inst_reg[11]_1 (\_T_2547[31]_i_4_n_0 ),
        .\wb_reg_inst_reg[22] (wb_reg_xcpt_i_2_n_0),
        .\wb_reg_inst_reg[7] (\wb_reg_inst_reg[7]_1 ),
        .\wb_reg_inst_reg[9] (\wb_reg_inst_reg[9]_3 ),
        .\wb_reg_inst_reg[9]_0 (\wb_reg_inst_reg[9]_0 ),
        .\wb_reg_inst_reg[9]_1 (\wb_reg_inst_reg[9]_1 ),
        .\wb_reg_inst_reg[9]_2 (\wb_reg_inst_reg[9]_2 ),
        .\wb_reg_inst_reg[9]_3 (\_T_2547[28]_i_3_n_0 ),
        .\wb_reg_inst_reg[9]_4 (\_T_2547[29]_i_3_n_0 ),
        .\wb_reg_inst_reg[9]_5 (\_T_2547[30]_i_3_n_0 ),
        .\wb_reg_inst_reg[9]_6 (\_T_2547[31]_i_5_n_0 ),
        .wb_reg_replay(wb_reg_replay),
        .wb_reg_replay_reg(wb_reg_replay_reg_2),
        .wb_reg_valid_reg(frontend_io_cpu_req_bits_speculative),
        .wb_reg_valid_reg_0(wb_reg_valid));
  FDRE #(
    .INIT(1'b0)) 
    \ex_cause_reg[0] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(csr_n_639),
        .Q(ex_cause[0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_cause_reg[1] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(csr_n_638),
        .Q(ex_cause[1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_cause_reg[2] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(csr_n_637),
        .Q(ex_cause[2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_cause_reg[3] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(csr_n_636),
        .Q(ex_cause[3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_cause_reg[63] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(csr_io_interrupt),
        .Q(ex_cause[63]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_ctrl_alu_dw_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ex_ctrl_alu_dw_reg_0),
        .Q(req_dw_reg),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_alu_fn_reg[0] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[3]_3 [0]),
        .Q(ex_ctrl_alu_fn[0]),
        .R(ibuf_n_50));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_alu_fn_reg[1] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[3]_3 [1]),
        .Q(ex_ctrl_alu_fn[1]),
        .R(ibuf_n_50));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_alu_fn_reg[2] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[3]_3 [2]),
        .Q(ex_ctrl_alu_fn[2]),
        .R(ibuf_n_50));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_alu_fn_reg[3] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[3]_3 [3]),
        .Q(Q),
        .R(ibuf_n_50));
  FDRE #(
    .INIT(1'b0)) 
    ex_ctrl_branch_reg
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[1]_1 ),
        .Q(ex_ctrl_branch),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_csr_reg[0] 
       (.C(host_clk),
        .CE(\<const1> ),
        .D(\ex_ctrl_csr_reg[0]_0 ),
        .Q(D[0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_csr_reg[1] 
       (.C(host_clk),
        .CE(\<const1> ),
        .D(\ex_ctrl_csr_reg[1]_0 ),
        .Q(D[1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_csr_reg[2] 
       (.C(host_clk),
        .CE(\<const1> ),
        .D(\ex_ctrl_csr_reg[2]_0 ),
        .Q(D[2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_ctrl_div_reg
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[1]_0 ),
        .Q(ex_ctrl_div),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_ctrl_fence_i_reg
       (.C(host_clk),
        .CE(_T_1790),
        .D(id_ctrl_fence_i),
        .Q(ex_ctrl_fence_i),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_ctrl_jal_reg
       (.C(host_clk),
        .CE(_T_1790),
        .D(id_ctrl_jal),
        .Q(ex_ctrl_jal),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_ctrl_jalr_reg
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[1] ),
        .Q(ex_ctrl_jalr),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_mem_cmd_reg[0] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[3]_1 [0]),
        .Q(\s1_req_cmd_reg[4] [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_mem_cmd_reg[1] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[3]_1 [1]),
        .Q(\s1_req_cmd_reg[4] [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_mem_cmd_reg[2] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[3]_1 [2]),
        .Q(\s1_req_cmd_reg[4] [2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_mem_cmd_reg[3] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[3]_1 [3]),
        .Q(\s1_req_cmd_reg[4] [3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_mem_cmd_reg[4] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(_T_1005[1]),
        .Q(\s1_req_cmd_reg[4] [4]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_ctrl_mem_reg
       (.C(host_clk),
        .CE(_T_1790),
        .D(id_ctrl_mem),
        .Q(ex_ctrl_mem),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_mem_type_reg[0] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[3]_2 [0]),
        .Q(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_mem_type_reg[1] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[3]_2 [1]),
        .Q(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_mem_type_reg[2] 
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ibuf_n_71),
        .Q(dcacheArb_io_requestor_1_req_bits_typ[2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_ctrl_rxs2_reg
       (.C(host_clk),
        .CE(_T_1790),
        .D(id_ctrl_rxs2),
        .Q(ex_ctrl_rxs2),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_sel_alu1_reg[0] 
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ibuf_n_74),
        .Q(\ex_ctrl_sel_alu1_reg[0]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_sel_alu1_reg[1] 
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ibuf_n_73),
        .Q(\ex_ctrl_sel_alu1_reg[1]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_sel_alu2_reg[0] 
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ibuf_n_72),
        .Q(ex_ctrl_sel_alu2[0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_sel_alu2_reg[1] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(buf__xcpt_pf_inst_reg_1),
        .Q(ex_ctrl_sel_alu2[1]),
        .R(ibuf_n_50));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_sel_imm_reg[0] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(nBufValid_reg_8[0]),
        .Q(\bypass_mux_1_reg[6]_1 [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_sel_imm_reg[1] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(nBufValid_reg_8[1]),
        .Q(\bypass_mux_1_reg[6]_1 [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_ctrl_sel_imm_reg[2] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(nBufValid_reg_8[2]),
        .Q(\bypass_mux_1_reg[6]_1 [2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_ctrl_wxd_reg
       (.C(host_clk),
        .CE(_T_1790),
        .D(id_ctrl_wxd),
        .Q(ex_ctrl_wxd),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_reg_flush_pipe_reg
       (.C(host_clk),
        .CE(_T_1790),
        .D(_T_1821),
        .Q(ex_reg_flush_pipe),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[10] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[3]),
        .Q(\mem_reg_inst_reg[31]_0 [3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[11] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[4]),
        .Q(\mem_reg_inst_reg[31]_0 [4]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[12] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_1142[0]),
        .Q(\ex_reg_inst_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[13] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_1142[1]),
        .Q(\ex_reg_inst_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[14] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_1031),
        .Q(\ex_reg_inst_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[15] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[5]),
        .Q(\ex_reg_inst_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[16] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[6]),
        .Q(\ex_reg_inst_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[17] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[7]),
        .Q(\ex_reg_inst_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[18] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[8]),
        .Q(\ex_reg_inst_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[19] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[9]),
        .Q(\ex_reg_inst_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[20] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[10]),
        .Q(_T_1710),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[21] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[11]),
        .Q(\ex_reg_inst_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[22] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[12]),
        .Q(\ex_reg_inst_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[23] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[13]),
        .Q(\ex_reg_inst_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[24] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[14]),
        .Q(\ex_reg_inst_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[25] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_877),
        .Q(\ex_reg_inst_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[26] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_909[0]),
        .Q(\mem_reg_inst_reg[31]_0 [5]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[27] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_909[1]),
        .Q(\mem_reg_inst_reg[31]_0 [6]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[28] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_909[2]),
        .Q(\ex_reg_inst_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[29] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_909[3]),
        .Q(\ex_reg_inst_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[30] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_1142[2]),
        .Q(\ex_reg_inst_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[31] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_909[4]),
        .Q(\mem_reg_inst_reg[31]_0 [7]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[7] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[0]),
        .Q(\mem_reg_inst_reg[31]_0 [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[8] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[1]),
        .Q(\mem_reg_inst_reg[31]_0 [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_inst_reg[9] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(_T_889[2]),
        .Q(\mem_reg_inst_reg[31]_0 [2]),
        .R(\<const0> ));
  LUT2 #(
    .INIT(4'h8)) 
    ex_reg_load_use_i_1
       (.I0(mem_ctrl_mem),
        .I1(ibuf_n_52),
        .O(id_load_use));
  FDRE #(
    .INIT(1'b0)) 
    ex_reg_load_use_reg
       (.C(host_clk),
        .CE(_T_1790),
        .D(id_load_use),
        .Q(ex_reg_load_use),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[10] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[10]),
        .Q(ex_reg_pc[10]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[11] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [3]),
        .Q(ex_reg_pc[11]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[12] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[12]),
        .Q(ex_reg_pc[12]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[13] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [4]),
        .Q(ex_reg_pc[13]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[14] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[14]),
        .Q(ex_reg_pc[14]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[15] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [5]),
        .Q(ex_reg_pc[15]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[16] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[16]),
        .Q(ex_reg_pc[16]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[17] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [6]),
        .Q(ex_reg_pc[17]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[18] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[18]),
        .Q(ex_reg_pc[18]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[19] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [7]),
        .Q(ex_reg_pc[19]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[1] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[1]),
        .Q(ex_reg_pc[1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[20] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[20]),
        .Q(ex_reg_pc[20]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[21] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [8]),
        .Q(ex_reg_pc[21]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[22] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[22]),
        .Q(ex_reg_pc[22]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[23] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [9]),
        .Q(ex_reg_pc[23]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[24] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[24]),
        .Q(ex_reg_pc[24]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[25] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [10]),
        .Q(ex_reg_pc[25]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[26] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[26]),
        .Q(ex_reg_pc[26]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[27] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [11]),
        .Q(ex_reg_pc[27]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[28] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[28]),
        .Q(ex_reg_pc[28]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[29] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [12]),
        .Q(ex_reg_pc[29]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[2] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[2]),
        .Q(ex_reg_pc[2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[30] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[30]),
        .Q(ex_reg_pc[30]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[31] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [13]),
        .Q(\mem_reg_pc_reg[31]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[32] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[32]),
        .Q(ex_reg_pc[32]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[33] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [14]),
        .Q(ex_reg_pc[33]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[34] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[34]),
        .Q(ex_reg_pc[34]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[35] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [15]),
        .Q(ex_reg_pc[35]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[36] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[36]),
        .Q(ex_reg_pc[36]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[37] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [16]),
        .Q(ex_reg_pc[37]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[38] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [17]),
        .Q(ex_reg_pc[38]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[39] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [18]),
        .Q(ex_reg_pc[39]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[3] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[3]),
        .Q(ex_reg_pc[3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[4] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[4]),
        .Q(ex_reg_pc[4]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[5] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [0]),
        .Q(ex_reg_pc[5]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[6] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[6]),
        .Q(ex_reg_pc[6]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[7] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [1]),
        .Q(ex_reg_pc[7]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[8] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(ibuf_io_pc[8]),
        .Q(ex_reg_pc[8]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_pc_reg[9] 
       (.C(host_clk),
        .CE(_T_1865),
        .D(\elts_0_pc_reg[39] [2]),
        .Q(ex_reg_pc[9]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_reg_replay_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ex_reg_replay0),
        .Q(ex_reg_replay),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_reg_rs_bypass_0_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ex_reg_rs_bypass_0_reg_1),
        .Q(ex_reg_rs_bypass_0_reg_0),
        .R(\<const0> ));
  LUT2 #(
    .INIT(4'h7)) 
    ex_reg_rs_bypass_1_i_1
       (.I0(ex_reg_rs_bypass_1_reg_0),
        .I1(ex_ctrl_wxd_reg_0),
        .O(_T_1844));
  FDRE #(
    .INIT(1'b0)) 
    ex_reg_rs_bypass_1_reg
       (.C(host_clk),
        .CE(_T_1790),
        .D(_T_1844),
        .Q(ex_reg_rs_bypass_1),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_lsb_0_reg[0] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[1]_3 [0]),
        .Q(ex_reg_rs_lsb_0[0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_lsb_0_reg[1] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(\buf__data_reg[1]_3 [1]),
        .Q(ex_reg_rs_lsb_0[1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_lsb_1_reg[0] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(ex_ctrl_wxd_reg_1[0]),
        .Q(\ex_reg_rs_lsb_1_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_lsb_1_reg[1] 
       (.C(host_clk),
        .CE(_T_1790),
        .D(ex_ctrl_wxd_reg_1[1]),
        .Q(\ex_reg_rs_lsb_1_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[0] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [0]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[10] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [10]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[11] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [11]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[12] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [12]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[13] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [13]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[14] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [14]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[15] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [15]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[16] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [16]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[17] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [17]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[18] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [18]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[19] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [19]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[1] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [1]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[20] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [20]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[21] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [21]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[22] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [22]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[23] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [23]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[24] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [24]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[25] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [25]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[26] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [26]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[27] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [27]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[28] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [28]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[29] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [29]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[2] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [2]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[30] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [30]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[30] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[31] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [31]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[31] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[32] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [32]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[32] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[33] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [33]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[33] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[34] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [34]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[34] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[35] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [35]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[35] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[36] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [36]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[36] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[37] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [37]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[37] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[38] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [38]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[38] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[39] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [39]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[39] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[3] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [3]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[40] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [40]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[40] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[41] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [41]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[41] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[42] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [42]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[42] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[43] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [43]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[43] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[44] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [44]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[44] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[45] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [45]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[45] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[46] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [46]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[46] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[47] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [47]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[47] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[48] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [48]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[48] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[49] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [49]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[49] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[4] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [4]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[50] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [50]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[50] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[51] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [51]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[51] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[52] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [52]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[52] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[53] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [53]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[53] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[54] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [54]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[54] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[55] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [55]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[55] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[56] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [56]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[56] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[57] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [57]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[57] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[58] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [58]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[58] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[59] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [59]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[59] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[5] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [5]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[60] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [60]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[60] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[61] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [61]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[61] ),
        .R(ex_reg_rs_bypass_0));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[6] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [6]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[7] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [7]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[8] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [8]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_0_reg[9] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_1 ),
        .D(\bypass_mux_2_reg[63]_2 [9]),
        .Q(\ex_reg_rs_msb_0_reg_n_0_[9] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[0] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[0]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[10] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[10]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[10] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[11] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[11]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[11] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[12] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[12]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[12] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[13] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[13]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[13] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[14] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[14]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[14] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[15] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[15]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[15] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[16] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[16]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[16] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[17] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[17]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[17] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[18] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[18]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[18] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[19] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[19]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[19] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[1] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[1]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[20] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[20]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[20] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[21] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[21]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[21] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[22] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[22]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[22] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[23] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[23]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[23] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[24] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[24]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[24] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[25] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[25]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[25] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[26] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[26]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[26] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[27] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[27]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[27] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[28] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[28]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[28] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[29] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[29]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[29] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[2] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[2]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[30] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[30]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[30] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[31] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[31]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[32] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[32]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[32] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[33] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[33]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[33] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[34] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[34]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[34] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[35] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[35]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[35] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[36] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[36]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[36] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[37] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[37]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[37] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[38] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[38]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[38] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[39] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[39]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[39] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[3] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[3]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[3] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[40] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[40]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[40] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[41] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[41]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[41] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[42] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[42]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[42] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[43] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[43]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[43] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[44] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[44]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[44] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[45] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[45]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[45] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[46] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[46]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[46] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[47] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[47]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[47] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[48] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[48]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[48] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[49] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[49]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[49] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[4] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[4]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[4] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[50] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[50]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[50] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[51] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[51]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[51] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[52] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[52]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[52] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[53] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[53]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[53] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[54] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[54]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[54] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[55] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[55]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[55] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[56] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[56]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[56] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[57] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[57]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[57] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[58] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[58]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[58] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[59] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[59]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[59] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[5] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[5]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[5] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[60] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[60]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[60] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[61] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[61]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[61] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[6] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[6]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[6] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[7] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[7]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[7] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[8] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[8]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[8] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \ex_reg_rs_msb_1_reg[9] 
       (.C(host_clk),
        .CE(\mem_reg_inst_reg[9]_0 ),
        .D(_T_1856[9]),
        .Q(\ex_reg_rs_msb_1_reg_n_0_[9] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_reg_rvc_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ex_reg_rvc_reg_1),
        .Q(mem_reg_rvc_reg_0),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_reg_valid_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(_T_1790),
        .Q(ex_reg_valid),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_reg_xcpt_interrupt_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ex_reg_xcpt_interrupt0),
        .Q(ex_reg_xcpt_interrupt),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    ex_reg_xcpt_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ibuf_n_50),
        .Q(ex_reg_xcpt),
        .R(\<const0> ));
  IBuf ibuf
       (.D({ibuf_io_pc[36],ibuf_io_pc[34],ibuf_io_pc[32],ibuf_io_pc[30],ibuf_io_pc[28],ibuf_io_pc[26],ibuf_io_pc[24],ibuf_io_pc[22],ibuf_io_pc[20],ibuf_io_pc[18],ibuf_io_pc[16],ibuf_io_pc[14],ibuf_io_pc[12],ibuf_io_pc[10],ibuf_io_pc[8],ibuf_io_pc[6],ibuf_io_pc[4:1]}),
        .E(_T_1865),
        .Q(\wb_reg_inst_reg[31]_0 [4:0]),
        .SR(ibuf_n_50),
        ._GEN_6(\bpu/_GEN_6 ),
        ._T_1031(_T_1031),
        ._T_134(_T_134),
        ._T_1573(_T_1573),
        .\_T_2547_reg[16] (\_T_2547_reg[16]_1 ),
        .\_T_2547_reg[31] ({_T_2549[31:17],\_T_2547_reg[16]_0 ,_T_2549[15:1]}),
        .\buf__data_reg[1]_0 (\buf__data_reg[1]_2 ),
        .\buf__data_reg[4]_0 (\buf__data_reg[4] ),
        .\buf__data_reg[4]_1 (\buf__data_reg[4]_0 ),
        .buf__pc(buf__pc),
        .buf__xcpt_ae_inst(buf__xcpt_ae_inst),
        .buf__xcpt_pf_inst_reg_0(buf__xcpt_pf_inst_reg),
        .buf__xcpt_pf_inst_reg_1(buf__xcpt_pf_inst_reg_2),
        .csr_io_bp_0_control_action(csr_io_bp_0_control_action),
        .dcacheArb_io_requestor_1_ordered(dcacheArb_io_requestor_1_ordered),
        .dcacheArb_io_requestor_1_req_bits_typ(dcacheArb_io_requestor_1_req_bits_typ[2]),
        .dcacheArb_io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),
        .dcache_blocked_reg(ex_ctrl_mem_reg_0),
        .\elts_0_data_reg[15] (\elts_0_data_reg[15] ),
        .\elts_0_pc_reg[37] (\elts_0_pc_reg[39] [16:0]),
        .elts_0_xcpt_ae_inst_reg(elts_0_xcpt_ae_inst_reg),
        .\ex_cause_reg[1] (\ex_cause_reg[1]_2 ),
        .\ex_cause_reg[1]_0 (\ex_cause_reg[1]_3 ),
        .\ex_cause_reg[1]_1 (\ex_cause_reg[1]_5 ),
        .\ex_cause_reg[1]_2 (\ex_cause_reg[1]_6 ),
        .\ex_cause_reg[1]_3 (\ex_cause_reg[1]_8 ),
        .\ex_cause_reg[1]_4 (\ex_cause_reg[1]_9 ),
        .\ex_cause_reg[1]_5 (\ex_cause_reg[1]_10 ),
        .\ex_cause_reg[1]_6 (\ex_cause_reg[1]_11 ),
        .\ex_cause_reg[1]_7 (\ex_cause_reg[1]_13 ),
        .\ex_cause_reg[1]_8 (\ex_cause_reg[1]_14 ),
        .\ex_cause_reg[1]_9 (\ex_cause_reg[1]_12 [1]),
        .\ex_cause_reg[2] (ibuf_n_65),
        .\ex_ctrl_csr_reg[2] (D),
        .ex_ctrl_div_reg(ex_ctrl_div),
        .ex_ctrl_jalr(ex_ctrl_jalr),
        .ex_ctrl_mem(ex_ctrl_mem),
        .ex_ctrl_mem_reg(_T_1790),
        .ex_ctrl_mem_reg_0(ex_ctrl_mem_reg_2),
        .ex_ctrl_mem_reg_1(ibuf_n_56),
        .ex_ctrl_mem_reg_10(ex_ctrl_mem_reg_10),
        .ex_ctrl_mem_reg_11(ibuf_n_68),
        .ex_ctrl_mem_reg_12(ex_ctrl_mem_reg_11),
        .ex_ctrl_mem_reg_2(ex_ctrl_mem_reg_3),
        .ex_ctrl_mem_reg_3(ex_ctrl_mem_reg_4),
        .ex_ctrl_mem_reg_4(ex_ctrl_mem_reg_5),
        .ex_ctrl_mem_reg_5(ex_ctrl_mem_reg_6),
        .ex_ctrl_mem_reg_6(ex_ctrl_mem_reg_7),
        .ex_ctrl_mem_reg_7(ex_ctrl_mem_reg_8),
        .ex_ctrl_mem_reg_8(ex_ctrl_mem_reg_9),
        .ex_ctrl_mem_reg_9(ibuf_n_64),
        .\ex_ctrl_mem_type_reg[2] (ibuf_n_71),
        .\ex_ctrl_sel_alu1_reg[0] (ibuf_n_74),
        .\ex_ctrl_sel_alu1_reg[0]_0 (\ex_ctrl_sel_alu1_reg[0]_0 ),
        .\ex_ctrl_sel_alu1_reg[1] (ibuf_n_73),
        .\ex_ctrl_sel_alu1_reg[1]_0 (\ex_ctrl_sel_alu1_reg[1]_0 ),
        .\ex_ctrl_sel_alu2_reg[0] (ibuf_n_72),
        .\ex_ctrl_sel_alu2_reg[0]_0 (ex_ctrl_sel_alu2[0]),
        .\ex_ctrl_sel_alu2_reg[1] (\ex_ctrl_sel_alu2_reg[1]_0 ),
        .\ex_ctrl_sel_alu2_reg[1]_0 (\ex_ctrl_sel_alu2_reg[1]_3 ),
        .ex_ctrl_wxd_reg(ex_ctrl_wxd),
        .\ex_reg_inst_reg[11] (\ex_reg_inst_reg[11]_0 ),
        .\ex_reg_inst_reg[11]_0 (\mem_reg_inst_reg[31]_0 [4:0]),
        .ex_reg_load_use_reg(ibuf_n_52),
        .\ex_reg_pc_reg[1] (_T_100),
        .\ex_reg_pc_reg[39] (\ex_reg_pc_reg[39]_0 ),
        .ex_reg_replay0(ex_reg_replay0),
        .ex_reg_replay_reg(buf__replay),
        .ex_reg_replay_reg_0(ibuf_n_47),
        .ex_reg_rs_bypass_1_reg(ex_reg_rs_bypass_1_reg_0),
        .\ex_reg_rs_lsb_0_reg[0] (\ex_reg_rs_lsb_0_reg[0]_0 ),
        .\ex_reg_rs_msb_0_reg[61] (ex_reg_rs_bypass_0),
        .ex_reg_valid_reg(ex_reg_valid),
        .frontend_io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
        .frontend_io_cpu_resp_bits_replay(frontend_io_cpu_resp_bits_replay),
        .frontend_io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),
        .frontend_io_cpu_resp_bits_xcpt_pf_inst(frontend_io_cpu_resp_bits_xcpt_pf_inst),
        .frontend_io_cpu_resp_valid(frontend_io_cpu_resp_valid),
        .host_clk(host_clk),
        .ibuf_io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
        .ibuf_io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
        .ibuf_io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
        .ibuf_io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
        .id_ctrl_sel_alu1(id_ctrl_sel_alu1),
        .id_reg_fence_reg(ibuf_n_70),
        .id_reg_fence_reg_0(div_n_368),
        .id_reg_fence_reg_1(id_reg_fence_reg_0),
        .\mem_ctrl_csr_reg[1] (mem_ctrl_csr[1:0]),
        .mem_ctrl_mem_reg(mem_ctrl_mem),
        .mem_ctrl_wxd(mem_ctrl_wxd),
        .\mem_reg_inst_reg[11] (\mem_reg_inst_reg[11]_0 ),
        .mem_reg_slow_bypass(mem_reg_slow_bypass),
        .mem_reg_valid_reg(mem_reg_replay_reg_0),
        .mem_reg_valid_reg_0(mem_reg_valid),
        .nBufValid_reg_0(nBufValid_reg),
        .nBufValid_reg_1(nBufValid_reg_2),
        .nBufValid_reg_2(nBufValid_reg_3),
        .nBufValid_reg_3(nBufValid_reg_4),
        .nBufValid_reg_4(nBufValid_reg_7),
        .nBufValid_reg_5(nBufValid_reg_9),
        .\reg_bp_0_address_reg[37] ({csr_io_bp_0_address,\reg_sscratch_reg[45] [3:2]}),
        .\reg_bp_0_control_tmatch_reg[1] (\ex_ctrl_sel_alu2_reg[1]_4 ),
        .\reg_misa_reg[12] (\reg_misa_reg[12]_0 ),
        .reg_mstatus_tvm_reg(reg_mstatus_tvm_reg),
        .reg_singleStepped_reg(csr_io_interrupt),
        .\s2_req_tag_reg[5] (\s2_req_tag_reg[5] ),
        .wb_ctrl_div(wb_ctrl_div),
        .wb_ctrl_mem_reg(wb_ctrl_mem),
        .wb_ctrl_wxd_reg(wb_ctrl_wxd),
        .\wb_reg_inst_reg[11] (\reg_bp_0_control_tmatch_reg[1] [4:0]),
        .\wb_reg_inst_reg[7] (\wb_reg_inst_reg[7]_0 ),
        .wb_reg_valid_reg(wb_reg_valid));
  FDRE #(
    .INIT(1'b0)) 
    id_reg_fence_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(ibuf_n_70),
        .Q(id_reg_fence_reg_0),
        .R(target_reset));
  LUT5 #(
    .INIT(32'hFF080000)) 
    invalidated_i_1
       (.I0(wb_ctrl_fence_i),
        .I1(wb_reg_valid),
        .I2(dcacheArb_io_requestor_1_s2_nack),
        .I3(invalidated),
        .I4(refill_valid),
        .O(invalidated_reg));
  LUT2 #(
    .INIT(4'h6)) 
    mem_br_taken__i_1
       (.I0(ex_ctrl_alu_fn[0]),
        .I1(\alu/_T_32 ),
        .O(alu_io_cmp_out));
  LUT6 #(
    .INIT(64'h8EB2FFFF8EB20000)) 
    mem_br_taken__i_2
       (.I0(\ex_reg_pc_reg[39]_1 ),
        .I1(alu_io_in2[62]),
        .I2(alu_io_in1[62]),
        .I3(ex_ctrl_alu_fn[1]),
        .I4(Q),
        .I5(\ex_ctrl_alu_fn_reg[3]_9 ),
        .O(\alu/_T_32 ));
  LUT3 #(
    .INIT(8'h69)) 
    mem_br_taken__i_5
       (.I0(Q),
        .I1(alu_io_in2[62]),
        .I2(alu_io_in1[62]),
        .O(mem_br_taken__reg_0));
  FDRE #(
    .INIT(1'b0)) 
    mem_br_taken__reg
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(alu_io_cmp_out),
        .Q(mem_br_taken_),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_ctrl_branch_reg
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_branch),
        .Q(mem_ctrl_branch),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_ctrl_csr_reg[0] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(D[0]),
        .Q(mem_ctrl_csr[0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_ctrl_csr_reg[1] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(D[1]),
        .Q(mem_ctrl_csr[1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_ctrl_csr_reg[2] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(D[2]),
        .Q(mem_ctrl_csr[2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_ctrl_div_reg
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_div),
        .Q(mem_ctrl_div),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_ctrl_fence_i_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(mem_ctrl_fence_i_reg_0),
        .Q(wb_ctrl_fence_i_reg_0),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_ctrl_jal_reg
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_jal),
        .Q(mem_ctrl_jal),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_ctrl_jalr_reg
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_jalr),
        .Q(mem_ctrl_jalr),
        .R(\<const0> ));
  LUT5 #(
    .INIT(32'h77777770)) 
    mem_ctrl_mem_i_1
       (.I0(mem_reg_flush_pipe),
        .I1(mem_reg_valid),
        .I2(ex_reg_xcpt_interrupt),
        .I3(ex_reg_valid),
        .I4(ex_reg_replay),
        .O(mem_ctrl_fp));
  FDRE #(
    .INIT(1'b0)) 
    mem_ctrl_mem_reg
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_mem),
        .Q(mem_ctrl_mem),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_ctrl_mem_type_reg[0] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .Q(\mem_ctrl_mem_type_reg_n_0_[0] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_ctrl_mem_type_reg[1] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .Q(\mem_ctrl_mem_type_reg_n_0_[1] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_ctrl_wxd_reg
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_ctrl_wxd),
        .Q(mem_ctrl_wxd),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_cause_reg[0] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_cause[0]),
        .Q(mem_reg_cause[0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_cause_reg[1] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_cause[1]),
        .Q(mem_reg_cause[1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_cause_reg[2] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_cause[2]),
        .Q(\wb_reg_cause_reg[3]_0 [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_cause_reg[3] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_cause[3]),
        .Q(\wb_reg_cause_reg[3]_0 [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_cause_reg[63] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_cause[63]),
        .Q(mem_reg_cause[63]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_reg_flush_pipe_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(mem_reg_flush_pipe_reg_0),
        .Q(mem_reg_flush_pipe),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[10] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\mem_reg_inst_reg[31]_0 [3]),
        .Q(\wb_reg_inst_reg[31]_0 [3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[11] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\mem_reg_inst_reg[31]_0 [4]),
        .Q(\wb_reg_inst_reg[31]_0 [4]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[12] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[12] ),
        .Q(\wb_reg_inst_reg[31]_0 [5]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[13] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[13] ),
        .Q(\wb_reg_inst_reg[31]_0 [6]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[14] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[14] ),
        .Q(\wb_reg_inst_reg[31]_0 [7]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[15] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[15] ),
        .Q(\wb_reg_inst_reg[31]_0 [8]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[16] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[16] ),
        .Q(\wb_reg_inst_reg[31]_0 [9]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[17] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[17] ),
        .Q(\wb_reg_inst_reg[31]_0 [10]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[18] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[18] ),
        .Q(\wb_reg_inst_reg[31]_0 [11]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[19] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[19] ),
        .Q(\wb_reg_inst_reg[31]_0 [12]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[20] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(_T_1710),
        .Q(\wb_reg_inst_reg[31]_0 [13]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[21] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[21] ),
        .Q(\wb_reg_inst_reg[31]_0 [14]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[22] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[22] ),
        .Q(\wb_reg_inst_reg[31]_0 [15]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[23] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[23] ),
        .Q(\wb_reg_inst_reg[31]_0 [16]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[24] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[24] ),
        .Q(\wb_reg_inst_reg[31]_0 [17]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[25] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[25] ),
        .Q(\wb_reg_inst_reg[31]_0 [18]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[26] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\mem_reg_inst_reg[31]_0 [5]),
        .Q(\wb_reg_inst_reg[31]_0 [19]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[27] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\mem_reg_inst_reg[31]_0 [6]),
        .Q(\wb_reg_inst_reg[31]_0 [20]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[28] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[28] ),
        .Q(\wb_reg_inst_reg[31]_0 [21]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[29] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[29] ),
        .Q(\wb_reg_inst_reg[31]_0 [22]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[30] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\ex_reg_inst_reg_n_0_[30] ),
        .Q(\wb_reg_inst_reg[31]_0 [23]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[31] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\mem_reg_inst_reg[31]_0 [7]),
        .Q(\wb_reg_inst_reg[31]_0 [24]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[7] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\mem_reg_inst_reg[31]_0 [0]),
        .Q(\wb_reg_inst_reg[31]_0 [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[8] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\mem_reg_inst_reg[31]_0 [1]),
        .Q(\wb_reg_inst_reg[31]_0 [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_inst_reg[9] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\mem_reg_inst_reg[31]_0 [2]),
        .Q(\wb_reg_inst_reg[31]_0 [2]),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h00000000F080F0B0)) 
    mem_reg_load_i_1
       (.I0(\s1_req_cmd_reg[4] [2]),
        .I1(\s1_req_cmd_reg[4] [1]),
        .I2(ex_ctrl_mem),
        .I3(\s1_req_cmd_reg[4] [3]),
        .I4(\s1_req_cmd_reg[4] [0]),
        .I5(\s1_req_cmd_reg[4] [4]),
        .O(_T_2269));
  FDRE #(
    .INIT(1'b0)) 
    mem_reg_load_reg
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(_T_2269),
        .Q(mem_reg_load),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[10] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[10]),
        .Q(\wb_reg_pc_reg[39]_0 [9]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[11] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[11]),
        .Q(\wb_reg_pc_reg[39]_0 [10]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[12] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[12]),
        .Q(\wb_reg_pc_reg[39]_0 [11]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[13] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[13]),
        .Q(\wb_reg_pc_reg[39]_0 [12]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[14] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[14]),
        .Q(\wb_reg_pc_reg[39]_0 [13]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[15] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[15]),
        .Q(\wb_reg_pc_reg[39]_0 [14]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[16] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[16]),
        .Q(\wb_reg_pc_reg[39]_0 [15]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[17] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[17]),
        .Q(\wb_reg_pc_reg[39]_0 [16]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[18] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[18]),
        .Q(\wb_reg_pc_reg[39]_0 [17]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[19] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[19]),
        .Q(\wb_reg_pc_reg[39]_0 [18]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[1] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[1]),
        .Q(\wb_reg_pc_reg[39]_0 [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[20] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[20]),
        .Q(\wb_reg_pc_reg[39]_0 [19]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[21] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[21]),
        .Q(\wb_reg_pc_reg[39]_0 [20]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[22] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[22]),
        .Q(\wb_reg_pc_reg[39]_0 [21]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[23] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[23]),
        .Q(\wb_reg_pc_reg[39]_0 [22]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[24] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[24]),
        .Q(\wb_reg_pc_reg[39]_0 [23]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[25] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[25]),
        .Q(\wb_reg_pc_reg[39]_0 [24]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[26] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[26]),
        .Q(\wb_reg_pc_reg[39]_0 [25]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[27] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[27]),
        .Q(\wb_reg_pc_reg[39]_0 [26]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[28] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[28]),
        .Q(\bypass_mux_2_reg[31]_0 [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[29] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[29]),
        .Q(\bypass_mux_2_reg[31]_0 [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[2] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[2]),
        .Q(\wb_reg_pc_reg[39]_0 [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[30] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[30]),
        .Q(\bypass_mux_2_reg[31]_0 [2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[31] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(\mem_reg_pc_reg[31]_0 ),
        .Q(\wb_reg_pc_reg[39]_0 [27]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[32] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[32]),
        .Q(\wb_reg_pc_reg[34]_0 [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[33] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[33]),
        .Q(\wb_reg_pc_reg[34]_0 [2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[34] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[34]),
        .Q(\wb_reg_pc_reg[34]_0 [3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[35] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[35]),
        .Q(\wb_reg_pc_reg[39]_0 [28]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[36] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[36]),
        .Q(\wb_reg_pc_reg[39]_0 [29]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[37] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[37]),
        .Q(\wb_reg_pc_reg[39]_0 [30]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[38] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[38]),
        .Q(\wb_reg_pc_reg[39]_0 [31]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[39] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[39]),
        .Q(\wb_reg_pc_reg[39]_0 [32]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[3] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[3]),
        .Q(\wb_reg_pc_reg[39]_0 [2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[4] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[4]),
        .Q(\wb_reg_pc_reg[39]_0 [3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[5] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[5]),
        .Q(\wb_reg_pc_reg[39]_0 [4]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[6] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[6]),
        .Q(\wb_reg_pc_reg[39]_0 [5]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[7] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[7]),
        .Q(\wb_reg_pc_reg[39]_0 [6]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[8] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[8]),
        .Q(\wb_reg_pc_reg[39]_0 [7]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_pc_reg[9] 
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(ex_reg_pc[9]),
        .Q(\wb_reg_pc_reg[39]_0 [8]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_reg_replay_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(mem_reg_replay0),
        .Q(mem_reg_replay),
        .R(\<const0> ));
  (* SOFT_HLUTNM = "soft_lutpair1823" *) 
  LUT4 #(
    .INIT(16'h02FE)) 
    \mem_reg_rs2[10]_i_1 
       (.I0(mem_reg_rs2[2]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(div_n_219),
        .O(mem_reg_rs20_in[10]));
  (* SOFT_HLUTNM = "soft_lutpair1824" *) 
  LUT4 #(
    .INIT(16'h333A)) 
    \mem_reg_rs2[11]_i_1 
       (.I0(mem_reg_rs2[3]),
        .I1(div_n_220),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .O(mem_reg_rs20_in[11]));
  (* SOFT_HLUTNM = "soft_lutpair1827" *) 
  LUT4 #(
    .INIT(16'h333A)) 
    \mem_reg_rs2[12]_i_1 
       (.I0(mem_reg_rs2[4]),
        .I1(div_n_221),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .O(mem_reg_rs20_in[12]));
  (* SOFT_HLUTNM = "soft_lutpair1828" *) 
  LUT4 #(
    .INIT(16'h333A)) 
    \mem_reg_rs2[13]_i_1 
       (.I0(mem_reg_rs2[5]),
        .I1(div_n_222),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .O(mem_reg_rs20_in[13]));
  (* SOFT_HLUTNM = "soft_lutpair1829" *) 
  LUT4 #(
    .INIT(16'h333A)) 
    \mem_reg_rs2[14]_i_1 
       (.I0(\divisor_reg[57] [1]),
        .I1(div_n_223),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .O(mem_reg_rs20_in[14]));
  (* SOFT_HLUTNM = "soft_lutpair1830" *) 
  LUT4 #(
    .INIT(16'h333A)) 
    \mem_reg_rs2[15]_i_1 
       (.I0(\divisor_reg[57] [2]),
        .I1(div_n_224),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .O(mem_reg_rs20_in[15]));
  (* SOFT_HLUTNM = "soft_lutpair1839" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mem_reg_rs2[16]_i_1 
       (.I0(mem_reg_rs2[16]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(mem_reg_rs2[0]),
        .O(mem_reg_rs20_in[16]));
  (* SOFT_HLUTNM = "soft_lutpair1838" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mem_reg_rs2[17]_i_1 
       (.I0(mem_reg_rs2[17]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(\divisor_reg[57] [0]),
        .O(mem_reg_rs20_in[17]));
  (* SOFT_HLUTNM = "soft_lutpair1837" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    \mem_reg_rs2[18]_i_1 
       (.I0(div_n_225),
        .I1(mem_reg_rs2[2]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .O(mem_reg_rs20_in[18]));
  (* SOFT_HLUTNM = "soft_lutpair1836" *) 
  LUT3 #(
    .INIT(8'h2E)) 
    \mem_reg_rs2[19]_i_1 
       (.I0(mem_reg_rs2[3]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(div_n_226),
        .O(mem_reg_rs20_in[19]));
  (* SOFT_HLUTNM = "soft_lutpair1835" *) 
  LUT3 #(
    .INIT(8'h2E)) 
    \mem_reg_rs2[20]_i_1 
       (.I0(mem_reg_rs2[4]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(div_n_227),
        .O(mem_reg_rs20_in[20]));
  (* SOFT_HLUTNM = "soft_lutpair1834" *) 
  LUT3 #(
    .INIT(8'h2E)) 
    \mem_reg_rs2[21]_i_1 
       (.I0(mem_reg_rs2[5]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(div_n_228),
        .O(mem_reg_rs20_in[21]));
  (* SOFT_HLUTNM = "soft_lutpair1833" *) 
  LUT3 #(
    .INIT(8'h2E)) 
    \mem_reg_rs2[22]_i_1 
       (.I0(\divisor_reg[57] [1]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(div_n_229),
        .O(mem_reg_rs20_in[22]));
  (* SOFT_HLUTNM = "soft_lutpair1831" *) 
  LUT3 #(
    .INIT(8'h2E)) 
    \mem_reg_rs2[23]_i_1 
       (.I0(\divisor_reg[57] [2]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(div_n_230),
        .O(mem_reg_rs20_in[23]));
  (* SOFT_HLUTNM = "soft_lutpair1825" *) 
  LUT5 #(
    .INIT(32'hFF3A003A)) 
    \mem_reg_rs2[24]_i_1 
       (.I0(mem_reg_rs2[0]),
        .I1(div_n_218),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[24]),
        .O(mem_reg_rs20_in[24]));
  (* SOFT_HLUTNM = "soft_lutpair1842" *) 
  LUT5 #(
    .INIT(32'hFF3A003A)) 
    \mem_reg_rs2[25]_i_1 
       (.I0(\divisor_reg[57] [0]),
        .I1(\mem_reg_rs2_reg[25]_0 ),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(\divisor_reg[57] [3]),
        .O(mem_reg_rs20_in[25]));
  (* SOFT_HLUTNM = "soft_lutpair1823" *) 
  LUT5 #(
    .INIT(32'hFF3A003A)) 
    \mem_reg_rs2[26]_i_1 
       (.I0(mem_reg_rs2[2]),
        .I1(div_n_219),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[26]),
        .O(mem_reg_rs20_in[26]));
  (* SOFT_HLUTNM = "soft_lutpair1824" *) 
  LUT5 #(
    .INIT(32'hFF3A003A)) 
    \mem_reg_rs2[27]_i_1 
       (.I0(mem_reg_rs2[3]),
        .I1(div_n_220),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[27]),
        .O(mem_reg_rs20_in[27]));
  (* SOFT_HLUTNM = "soft_lutpair1827" *) 
  LUT5 #(
    .INIT(32'hFF3A003A)) 
    \mem_reg_rs2[28]_i_1 
       (.I0(mem_reg_rs2[4]),
        .I1(div_n_221),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[28]),
        .O(mem_reg_rs20_in[28]));
  (* SOFT_HLUTNM = "soft_lutpair1828" *) 
  LUT5 #(
    .INIT(32'hFF3A003A)) 
    \mem_reg_rs2[29]_i_1 
       (.I0(mem_reg_rs2[5]),
        .I1(div_n_222),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[29]),
        .O(mem_reg_rs20_in[29]));
  (* SOFT_HLUTNM = "soft_lutpair1829" *) 
  LUT5 #(
    .INIT(32'hFF3A003A)) 
    \mem_reg_rs2[30]_i_1 
       (.I0(\divisor_reg[57] [1]),
        .I1(div_n_223),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[30]),
        .O(mem_reg_rs20_in[30]));
  (* SOFT_HLUTNM = "soft_lutpair1830" *) 
  LUT5 #(
    .INIT(32'hFF3A003A)) 
    \mem_reg_rs2[31]_i_1 
       (.I0(\divisor_reg[57] [2]),
        .I1(div_n_224),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[31]),
        .O(mem_reg_rs20_in[31]));
  LUT4 #(
    .INIT(16'hEA2A)) 
    \mem_reg_rs2[32]_i_1 
       (.I0(mem_reg_rs2[0]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[32]),
        .O(mem_reg_rs20_in[32]));
  LUT4 #(
    .INIT(16'hEA2A)) 
    \mem_reg_rs2[33]_i_1 
       (.I0(\divisor_reg[57] [0]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[33]),
        .O(mem_reg_rs20_in[33]));
  LUT4 #(
    .INIT(16'hEA2A)) 
    \mem_reg_rs2[34]_i_1 
       (.I0(mem_reg_rs2[2]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[34]),
        .O(mem_reg_rs20_in[34]));
  LUT4 #(
    .INIT(16'hEA2A)) 
    \mem_reg_rs2[35]_i_1 
       (.I0(mem_reg_rs2[3]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[35]),
        .O(mem_reg_rs20_in[35]));
  LUT4 #(
    .INIT(16'hEA2A)) 
    \mem_reg_rs2[36]_i_1 
       (.I0(mem_reg_rs2[4]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[36]),
        .O(mem_reg_rs20_in[36]));
  LUT4 #(
    .INIT(16'hEA2A)) 
    \mem_reg_rs2[37]_i_1 
       (.I0(mem_reg_rs2[5]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[37]),
        .O(mem_reg_rs20_in[37]));
  LUT4 #(
    .INIT(16'hEA2A)) 
    \mem_reg_rs2[38]_i_1 
       (.I0(\divisor_reg[57] [1]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[38]),
        .O(mem_reg_rs20_in[38]));
  LUT4 #(
    .INIT(16'hEA2A)) 
    \mem_reg_rs2[39]_i_1 
       (.I0(\divisor_reg[57] [2]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[39]),
        .O(mem_reg_rs20_in[39]));
  LUT5 #(
    .INIT(32'hC00ACFFA)) 
    \mem_reg_rs2[40]_i_1 
       (.I0(mem_reg_rs2[0]),
        .I1(mem_reg_rs2[40]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(div_n_218),
        .O(mem_reg_rs20_in[40]));
  LUT5 #(
    .INIT(32'hC00ACFFA)) 
    \mem_reg_rs2[42]_i_1 
       (.I0(mem_reg_rs2[2]),
        .I1(mem_reg_rs2[42]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(div_n_219),
        .O(mem_reg_rs20_in[42]));
  LUT5 #(
    .INIT(32'hC55FC550)) 
    \mem_reg_rs2[43]_i_1 
       (.I0(div_n_220),
        .I1(mem_reg_rs2[43]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[3]),
        .O(mem_reg_rs20_in[43]));
  LUT5 #(
    .INIT(32'hC55FC550)) 
    \mem_reg_rs2[44]_i_1 
       (.I0(div_n_221),
        .I1(mem_reg_rs2[44]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[4]),
        .O(mem_reg_rs20_in[44]));
  LUT5 #(
    .INIT(32'hC55FC550)) 
    \mem_reg_rs2[45]_i_1 
       (.I0(div_n_222),
        .I1(mem_reg_rs2[45]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[5]),
        .O(mem_reg_rs20_in[45]));
  LUT5 #(
    .INIT(32'hC55FC550)) 
    \mem_reg_rs2[46]_i_1 
       (.I0(div_n_223),
        .I1(mem_reg_rs2[46]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(\divisor_reg[57] [1]),
        .O(mem_reg_rs20_in[46]));
  LUT5 #(
    .INIT(32'hC55FC550)) 
    \mem_reg_rs2[47]_i_1 
       (.I0(div_n_224),
        .I1(mem_reg_rs2[47]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(\divisor_reg[57] [2]),
        .O(mem_reg_rs20_in[47]));
  (* SOFT_HLUTNM = "soft_lutpair1839" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mem_reg_rs2[48]_i_1 
       (.I0(mem_reg_rs2[48]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I2(mem_reg_rs2[16]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(mem_reg_rs2[0]),
        .O(mem_reg_rs20_in[48]));
  (* SOFT_HLUTNM = "soft_lutpair1838" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \mem_reg_rs2[49]_i_1 
       (.I0(mem_reg_rs2[49]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I2(mem_reg_rs2[17]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(\divisor_reg[57] [0]),
        .O(mem_reg_rs20_in[49]));
  (* SOFT_HLUTNM = "soft_lutpair1837" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    \mem_reg_rs2[50]_i_1 
       (.I0(div_n_234),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I2(div_n_225),
        .I3(mem_reg_rs2[2]),
        .I4(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .O(mem_reg_rs20_in[50]));
  (* SOFT_HLUTNM = "soft_lutpair1836" *) 
  LUT5 #(
    .INIT(32'h30AA3FAA)) 
    \mem_reg_rs2[51]_i_1 
       (.I0(mem_reg_rs2[3]),
        .I1(div_n_235),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(div_n_226),
        .O(mem_reg_rs20_in[51]));
  (* SOFT_HLUTNM = "soft_lutpair1835" *) 
  LUT5 #(
    .INIT(32'h30AA3FAA)) 
    \mem_reg_rs2[52]_i_1 
       (.I0(mem_reg_rs2[4]),
        .I1(div_n_236),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(div_n_227),
        .O(mem_reg_rs20_in[52]));
  (* SOFT_HLUTNM = "soft_lutpair1834" *) 
  LUT5 #(
    .INIT(32'h30AA3FAA)) 
    \mem_reg_rs2[53]_i_1 
       (.I0(mem_reg_rs2[5]),
        .I1(div_n_237),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(div_n_228),
        .O(mem_reg_rs20_in[53]));
  (* SOFT_HLUTNM = "soft_lutpair1833" *) 
  LUT5 #(
    .INIT(32'h30AA3FAA)) 
    \mem_reg_rs2[54]_i_1 
       (.I0(\divisor_reg[57] [1]),
        .I1(div_n_238),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(div_n_229),
        .O(mem_reg_rs20_in[54]));
  (* SOFT_HLUTNM = "soft_lutpair1831" *) 
  LUT5 #(
    .INIT(32'h30AA3FAA)) 
    \mem_reg_rs2[55]_i_1 
       (.I0(\divisor_reg[57] [2]),
        .I1(div_n_239),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I4(div_n_230),
        .O(mem_reg_rs20_in[55]));
  LUT6 #(
    .INIT(64'hF0AA00CCF0AAFFCC)) 
    \mem_reg_rs2[56]_i_1 
       (.I0(mem_reg_rs2[24]),
        .I1(mem_reg_rs2[0]),
        .I2(mem_reg_rs2[56]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I4(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I5(div_n_218),
        .O(mem_reg_rs20_in[56]));
  LUT6 #(
    .INIT(64'hF0AA00CCF0AAFFCC)) 
    \mem_reg_rs2[58]_i_1 
       (.I0(mem_reg_rs2[26]),
        .I1(mem_reg_rs2[2]),
        .I2(mem_reg_rs2[58]),
        .I3(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I4(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I5(div_n_219),
        .O(mem_reg_rs20_in[58]));
  LUT6 #(
    .INIT(64'hAFAFA0A03F303F30)) 
    \mem_reg_rs2[59]_i_1 
       (.I0(mem_reg_rs2[59]),
        .I1(div_n_220),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[3]),
        .I4(mem_reg_rs2[27]),
        .I5(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .O(mem_reg_rs20_in[59]));
  LUT6 #(
    .INIT(64'hAFAFA0A03F303F30)) 
    \mem_reg_rs2[60]_i_1 
       (.I0(mem_reg_rs2[60]),
        .I1(div_n_221),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[4]),
        .I4(mem_reg_rs2[28]),
        .I5(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .O(mem_reg_rs20_in[60]));
  LUT6 #(
    .INIT(64'hAFAFA0A03F303F30)) 
    \mem_reg_rs2[61]_i_1 
       (.I0(mem_reg_rs2[61]),
        .I1(div_n_222),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(mem_reg_rs2[5]),
        .I4(mem_reg_rs2[29]),
        .I5(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .O(mem_reg_rs20_in[61]));
  LUT6 #(
    .INIT(64'hAFAFA0A03F303F30)) 
    \mem_reg_rs2[62]_i_1 
       (.I0(mem_reg_rs2[62]),
        .I1(div_n_223),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(\divisor_reg[57] [1]),
        .I4(mem_reg_rs2[30]),
        .I5(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .O(mem_reg_rs20_in[62]));
  LUT3 #(
    .INIT(8'h80)) 
    \mem_reg_rs2[63]_i_1 
       (.I0(mem_ctrl_fp),
        .I1(ex_ctrl_rxs2),
        .I2(ex_ctrl_mem),
        .O(\mem_reg_rs2[63]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFA0A03F303F30)) 
    \mem_reg_rs2[63]_i_2 
       (.I0(mem_reg_rs2[63]),
        .I1(div_n_224),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(\divisor_reg[57] [2]),
        .I4(mem_reg_rs2[31]),
        .I5(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .O(mem_reg_rs20_in[63]));
  (* SOFT_HLUTNM = "soft_lutpair1825" *) 
  LUT4 #(
    .INIT(16'h02FE)) 
    \mem_reg_rs2[8]_i_1 
       (.I0(mem_reg_rs2[0]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(div_n_218),
        .O(mem_reg_rs20_in[8]));
  (* SOFT_HLUTNM = "soft_lutpair1842" *) 
  LUT4 #(
    .INIT(16'h02FE)) 
    \mem_reg_rs2[9]_i_1 
       (.I0(\divisor_reg[57] [0]),
        .I1(dcacheArb_io_requestor_1_req_bits_typ[1]),
        .I2(dcacheArb_io_requestor_1_req_bits_typ[0]),
        .I3(\mem_reg_rs2_reg[25]_0 ),
        .O(mem_reg_rs20_in[9]));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[0] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs2[0]),
        .Q(\a_data_reg[63] [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[10] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[10]),
        .Q(\a_data_reg[63] [10]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[11] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[11]),
        .Q(\a_data_reg[63] [11]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[12] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[12]),
        .Q(\a_data_reg[63] [12]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[13] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[13]),
        .Q(\a_data_reg[63] [13]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[14] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[14]),
        .Q(\a_data_reg[63] [14]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[15] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[15]),
        .Q(\a_data_reg[63] [15]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[16] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[16]),
        .Q(\a_data_reg[63] [16]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[17] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[17]),
        .Q(\a_data_reg[63] [17]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[18] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[18]),
        .Q(\a_data_reg[63] [18]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[19] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[19]),
        .Q(\a_data_reg[63] [19]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[1] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(\divisor_reg[57] [0]),
        .Q(\a_data_reg[63] [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[20] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[20]),
        .Q(\a_data_reg[63] [20]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[21] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[21]),
        .Q(\a_data_reg[63] [21]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[22] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[22]),
        .Q(\a_data_reg[63] [22]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[23] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[23]),
        .Q(\a_data_reg[63] [23]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[24] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[24]),
        .Q(\a_data_reg[63] [24]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[25] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[25]),
        .Q(\a_data_reg[63] [25]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[26] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[26]),
        .Q(\a_data_reg[63] [26]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[27] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[27]),
        .Q(\a_data_reg[63] [27]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[28] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[28]),
        .Q(\a_data_reg[63] [28]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[29] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[29]),
        .Q(\a_data_reg[63] [29]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[2] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs2[2]),
        .Q(\a_data_reg[63] [2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[30] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[30]),
        .Q(\a_data_reg[63] [30]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[31] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[31]),
        .Q(\a_data_reg[63] [31]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[32] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[32]),
        .Q(\a_data_reg[63] [32]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[33] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[33]),
        .Q(\a_data_reg[63] [33]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[34] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[34]),
        .Q(\a_data_reg[63] [34]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[35] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[35]),
        .Q(\a_data_reg[63] [35]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[36] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[36]),
        .Q(\a_data_reg[63] [36]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[37] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[37]),
        .Q(\a_data_reg[63] [37]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[38] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[38]),
        .Q(\a_data_reg[63] [38]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[39] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[39]),
        .Q(\a_data_reg[63] [39]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[3] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs2[3]),
        .Q(\a_data_reg[63] [3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[40] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[40]),
        .Q(\a_data_reg[63] [40]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[41] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(\ex_ctrl_mem_type_reg[0]_0 [0]),
        .Q(\a_data_reg[63] [41]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[42] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[42]),
        .Q(\a_data_reg[63] [42]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[43] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[43]),
        .Q(\a_data_reg[63] [43]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[44] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[44]),
        .Q(\a_data_reg[63] [44]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[45] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[45]),
        .Q(\a_data_reg[63] [45]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[46] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[46]),
        .Q(\a_data_reg[63] [46]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[47] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[47]),
        .Q(\a_data_reg[63] [47]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[48] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[48]),
        .Q(\a_data_reg[63] [48]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[49] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[49]),
        .Q(\a_data_reg[63] [49]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[4] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs2[4]),
        .Q(\a_data_reg[63] [4]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[50] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[50]),
        .Q(\a_data_reg[63] [50]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[51] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[51]),
        .Q(\a_data_reg[63] [51]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[52] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[52]),
        .Q(\a_data_reg[63] [52]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[53] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[53]),
        .Q(\a_data_reg[63] [53]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[54] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[54]),
        .Q(\a_data_reg[63] [54]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[55] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[55]),
        .Q(\a_data_reg[63] [55]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[56] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[56]),
        .Q(\a_data_reg[63] [56]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[57] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(\ex_ctrl_mem_type_reg[0]_0 [1]),
        .Q(\a_data_reg[63] [57]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[58] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[58]),
        .Q(\a_data_reg[63] [58]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[59] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[59]),
        .Q(\a_data_reg[63] [59]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[5] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs2[5]),
        .Q(\a_data_reg[63] [5]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[60] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[60]),
        .Q(\a_data_reg[63] [60]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[61] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[61]),
        .Q(\a_data_reg[63] [61]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[62] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[62]),
        .Q(\a_data_reg[63] [62]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[63] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[63]),
        .Q(\a_data_reg[63] [63]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[6] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(\divisor_reg[57] [1]),
        .Q(\a_data_reg[63] [6]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[7] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(\divisor_reg[57] [2]),
        .Q(\a_data_reg[63] [7]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[8] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[8]),
        .Q(\a_data_reg[63] [8]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \mem_reg_rs2_reg[9] 
       (.C(host_clk),
        .CE(\mem_reg_rs2[63]_i_1_n_0 ),
        .D(mem_reg_rs20_in[9]),
        .Q(\a_data_reg[63] [9]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_reg_rvc_reg
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(mem_reg_rvc_reg_0),
        .Q(mem_reg_rvc),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_reg_sfence_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(mem_reg_sfence_reg_1),
        .Q(mem_reg_sfence),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_reg_slow_bypass_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(mem_reg_slow_bypass_reg_1),
        .Q(mem_reg_slow_bypass),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h44444444400C0400)) 
    mem_reg_store_i_1
       (.I0(\s1_req_cmd_reg[4] [4]),
        .I1(ex_ctrl_mem),
        .I2(\s1_req_cmd_reg[4] [1]),
        .I3(\s1_req_cmd_reg[4] [2]),
        .I4(\s1_req_cmd_reg[4] [0]),
        .I5(\s1_req_cmd_reg[4] [3]),
        .O(_T_2305));
  FDRE #(
    .INIT(1'b0)) 
    mem_reg_store_reg
       (.C(host_clk),
        .CE(mem_ctrl_fp),
        .D(_T_2305),
        .Q(mem_reg_store),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_reg_valid_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(_T_2222),
        .Q(mem_reg_valid),
        .R(\<const0> ));
  (* SOFT_HLUTNM = "soft_lutpair1884" *) 
  LUT2 #(
    .INIT(4'h2)) 
    mem_reg_xcpt_interrupt_i_1
       (.I0(ex_reg_xcpt_interrupt),
        .I1(mem_reg_replay_reg_0),
        .O(mem_reg_xcpt_interrupt0));
  FDRE #(
    .INIT(1'b0)) 
    mem_reg_xcpt_interrupt_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(mem_reg_xcpt_interrupt0),
        .Q(mem_reg_xcpt_interrupt),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    mem_reg_xcpt_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(mem_reg_xcpt0),
        .Q(mem_reg_xcpt),
        .R(\<const0> ));
  (* SOFT_HLUTNM = "soft_lutpair1821" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \reg_sptbr_ppn[19]_i_4 
       (.I0(\reg_bp_0_control_tmatch_reg[1] [7]),
        .I1(\reg_bp_0_control_tmatch_reg[1] [5]),
        .I2(\reg_bp_0_control_tmatch_reg[1] [6]),
        .O(\reg_sptbr_ppn[19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[10]_i_4 
       (.I0(p_0_in[10]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[10] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [9]),
        .O(\s1_pc[10]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[11]_i_4 
       (.I0(p_0_in[11]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[11] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [10]),
        .O(\s1_pc[11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[12]_i_5 
       (.I0(p_0_in[12]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[12] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [11]),
        .O(\s1_pc[12]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[13]_i_4 
       (.I0(p_0_in[13]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[13] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [12]),
        .O(\s1_pc[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[14]_i_4 
       (.I0(p_0_in[14]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[14] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [13]),
        .O(\s1_pc[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[15]_i_4 
       (.I0(p_0_in[15]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[15] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [14]),
        .O(\s1_pc[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[16]_i_5 
       (.I0(p_0_in[16]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[16] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [15]),
        .O(\s1_pc[16]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[17]_i_4 
       (.I0(p_0_in[17]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[17] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [16]),
        .O(\s1_pc[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[18]_i_4 
       (.I0(p_0_in[18]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[18] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [17]),
        .O(\s1_pc[18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[19]_i_4 
       (.I0(p_0_in[19]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[19] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [18]),
        .O(\s1_pc[19]_i_4_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1862" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \s1_pc[1]_i_3 
       (.I0(p_0_in[1]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\mem_reg_rs2_reg[3]_1 [0]),
        .O(\s1_pc[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[20]_i_5 
       (.I0(p_0_in[20]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[20] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [19]),
        .O(\s1_pc[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[21]_i_4 
       (.I0(p_0_in[21]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[21] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [20]),
        .O(\s1_pc[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[22]_i_4 
       (.I0(p_0_in[22]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[22] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [21]),
        .O(\s1_pc[22]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[23]_i_4 
       (.I0(p_0_in[23]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[23] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [22]),
        .O(\s1_pc[23]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[24]_i_5 
       (.I0(p_0_in[24]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[24] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [23]),
        .O(\s1_pc[24]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[25]_i_4 
       (.I0(p_0_in[25]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[25] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [24]),
        .O(\s1_pc[25]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[26]_i_4 
       (.I0(p_0_in[26]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[26] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [25]),
        .O(\s1_pc[26]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[27]_i_4 
       (.I0(p_0_in[27]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[27] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [26]),
        .O(\s1_pc[27]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[28]_i_5 
       (.I0(p_0_in[28]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[28] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [27]),
        .O(\s1_pc[28]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[29]_i_4 
       (.I0(p_0_in[29]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[29] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [28]),
        .O(\s1_pc[29]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[2]_i_4 
       (.I0(p_0_in[2]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[2] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [1]),
        .O(\s1_pc[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[30]_i_4 
       (.I0(p_0_in[30]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[30] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [29]),
        .O(\s1_pc[30]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[31]_i_4 
       (.I0(p_0_in[31]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[31] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [30]),
        .O(\s1_pc[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[32]_i_4 
       (.I0(p_0_in[32]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[32] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [31]),
        .O(\s1_pc[32]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[33]_i_3 
       (.I0(p_0_in[33]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[33] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [32]),
        .O(\s1_pc[33]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[34]_i_3 
       (.I0(p_0_in[34]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[34] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [33]),
        .O(\s1_pc[34]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[35]_i_3 
       (.I0(p_0_in[35]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[35] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [34]),
        .O(\s1_pc[35]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[36]_i_4 
       (.I0(p_0_in[36]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[36] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [35]),
        .O(\s1_pc[36]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[37]_i_3 
       (.I0(p_0_in[37]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[37] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [36]),
        .O(\s1_pc[37]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[38]_i_3 
       (.I0(p_0_in[38]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_2_reg[38]_0 ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [37]),
        .O(\s1_pc[38]_i_3_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \s1_pc[39]_i_15 
       (.I0(_T_2177[24]),
        .O(\s1_pc_reg[39]_5 ));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_pc[39]_i_17 
       (.I0(_T_2177[21]),
        .I1(_T_2177[22]),
        .I2(_T_2177[23]),
        .O(\s1_pc_reg[39]_2 [3]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_pc[39]_i_18 
       (.I0(_T_2177[18]),
        .I1(_T_2177[19]),
        .I2(_T_2177[20]),
        .O(\s1_pc_reg[39]_2 [2]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_pc[39]_i_19 
       (.I0(_T_2177[15]),
        .I1(_T_2177[16]),
        .I2(_T_2177[17]),
        .O(\s1_pc_reg[39]_2 [1]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_pc[39]_i_20 
       (.I0(_T_2177[12]),
        .I1(_T_2177[13]),
        .I2(_T_2177[14]),
        .O(\s1_pc_reg[39]_2 [0]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_pc[39]_i_22 
       (.I0(_T_2177[22]),
        .I1(_T_2177[23]),
        .I2(_T_2177[21]),
        .O(\s1_pc_reg[39]_4 [3]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_pc[39]_i_23 
       (.I0(_T_2177[19]),
        .I1(_T_2177[20]),
        .I2(_T_2177[18]),
        .O(\s1_pc_reg[39]_4 [2]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_pc[39]_i_24 
       (.I0(_T_2177[16]),
        .I1(_T_2177[17]),
        .I2(_T_2177[15]),
        .O(\s1_pc_reg[39]_4 [1]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_pc[39]_i_25 
       (.I0(_T_2177[13]),
        .I1(_T_2177[14]),
        .I2(_T_2177[12]),
        .O(\s1_pc_reg[39]_4 [0]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_pc[39]_i_26 
       (.I0(_T_2177[9]),
        .I1(_T_2177[10]),
        .I2(_T_2177[11]),
        .O(\s1_pc_reg[39]_1 [3]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_pc[39]_i_27 
       (.I0(_T_2177[6]),
        .I1(_T_2177[7]),
        .I2(_T_2177[8]),
        .O(\s1_pc_reg[39]_1 [2]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_pc[39]_i_28 
       (.I0(_T_2177[3]),
        .I1(_T_2177[4]),
        .I2(_T_2177[5]),
        .O(\s1_pc_reg[39]_1 [1]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_pc[39]_i_29 
       (.I0(_T_2177[0]),
        .I1(_T_2177[1]),
        .I2(_T_2177[2]),
        .O(\s1_pc_reg[39]_1 [0]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_pc[39]_i_30 
       (.I0(_T_2177[10]),
        .I1(_T_2177[11]),
        .I2(_T_2177[9]),
        .O(\s1_pc_reg[39]_3 [3]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_pc[39]_i_31 
       (.I0(_T_2177[7]),
        .I1(_T_2177[8]),
        .I2(_T_2177[6]),
        .O(\s1_pc_reg[39]_3 [2]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_pc[39]_i_32 
       (.I0(_T_2177[4]),
        .I1(_T_2177[5]),
        .I2(_T_2177[3]),
        .O(\s1_pc_reg[39]_3 [1]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_pc[39]_i_33 
       (.I0(_T_2177[1]),
        .I1(_T_2177[2]),
        .I2(_T_2177[0]),
        .O(\s1_pc_reg[39]_3 [0]));
  LUT6 #(
    .INIT(64'hB8B8B888B8B8B8BB)) 
    \s1_pc[39]_i_4 
       (.I0(p_0_in[39]),
        .I1(core__707_i_3_n_0),
        .I2(_T_2177[0]),
        .I3(\bypass_mux_1_reg[63]_1 ),
        .I4(\bypass_mux_1_reg[63]_2 ),
        .I5(\bypass_mux_2_reg[38]_0 ),
        .O(\s1_pc[39]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[3]_i_4 
       (.I0(p_0_in[3]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\mem_reg_rs2_reg[3]_1 [1]),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [2]),
        .O(\s1_pc[3]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \s1_pc[3]_i_7 
       (.I0(wb_reg_valid),
        .I1(\reg_sscratch_reg[59] [2]),
        .I2(\reg_sscratch_reg[59] [1]),
        .I3(\reg_sscratch_reg[59] [0]),
        .I4(\reg_sptbr_ppn[19]_i_4_n_0 ),
        .O(\s1_pc[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[4]_i_4 
       (.I0(p_0_in[4]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[4] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [3]),
        .O(\s1_pc[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[5]_i_3 
       (.I0(p_0_in[5]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[5] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [4]),
        .O(\s1_pc[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[6]_i_4 
       (.I0(p_0_in[6]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[6] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [5]),
        .O(\s1_pc[6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[7]_i_4 
       (.I0(p_0_in[7]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[7] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [6]),
        .O(\s1_pc[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[8]_i_5 
       (.I0(p_0_in[8]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[8] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [7]),
        .O(\s1_pc[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFE02FFFFFE020000)) 
    \s1_pc[9]_i_4 
       (.I0(p_0_in[9]),
        .I1(mem_reg_sfence),
        .I2(mem_ctrl_jalr),
        .I3(\bypass_mux_1_reg_n_0_[9] ),
        .I4(wb_reg_replay_reg_1),
        .I5(\reg_dpc_reg[39] [8]),
        .O(\s1_pc[9]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_req_addr[39]_i_10 
       (.I0(\s1_req_addr_reg[39] [13]),
        .I1(\s1_req_addr_reg[39] [14]),
        .I2(_T_2770[20]),
        .O(\s1_req_addr_reg[39]_2 [2]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_req_addr[39]_i_11 
       (.I0(\s1_req_addr_reg[39] [11]),
        .I1(\s1_req_addr_reg[39] [12]),
        .I2(_T_2770[17]),
        .O(\s1_req_addr_reg[39]_2 [1]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_req_addr[39]_i_12 
       (.I0(\s1_req_addr_reg[39] [9]),
        .I1(\s1_req_addr_reg[39] [10]),
        .I2(_T_2770[14]),
        .O(\s1_req_addr_reg[39]_2 [0]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_req_addr[39]_i_14 
       (.I0(\s1_req_addr_reg[39] [15]),
        .I1(\s1_req_addr_reg[39] [16]),
        .I2(\s1_req_addr_reg[39] [17]),
        .O(\s1_req_addr_reg[39]_3 [3]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_req_addr[39]_i_15 
       (.I0(\s1_req_addr_reg[39] [13]),
        .I1(\s1_req_addr_reg[39] [14]),
        .I2(_T_2770[20]),
        .O(\s1_req_addr_reg[39]_3 [2]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_req_addr[39]_i_16 
       (.I0(\s1_req_addr_reg[39] [11]),
        .I1(\s1_req_addr_reg[39] [12]),
        .I2(_T_2770[17]),
        .O(\s1_req_addr_reg[39]_3 [1]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_req_addr[39]_i_17 
       (.I0(\s1_req_addr_reg[39] [9]),
        .I1(\s1_req_addr_reg[39] [10]),
        .I2(_T_2770[14]),
        .O(\s1_req_addr_reg[39]_3 [0]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_req_addr[39]_i_18 
       (.I0(_T_2770[9]),
        .I1(\s1_req_addr_reg[39] [7]),
        .I2(\s1_req_addr_reg[39] [8]),
        .O(\s1_req_addr_reg[39]_0 [3]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_req_addr[39]_i_19 
       (.I0(_T_2770[6]),
        .I1(\s1_req_addr_reg[39] [5]),
        .I2(\s1_req_addr_reg[39] [6]),
        .O(\s1_req_addr_reg[39]_0 [2]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_req_addr[39]_i_20 
       (.I0(\s1_req_addr_reg[39] [2]),
        .I1(\s1_req_addr_reg[39] [3]),
        .I2(\s1_req_addr_reg[39] [4]),
        .O(\s1_req_addr_reg[39]_0 [1]));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_req_addr[39]_i_21 
       (.I0(\s1_req_addr_reg[39] [0]),
        .I1(_T_2770[1]),
        .I2(\s1_req_addr_reg[39] [1]),
        .O(\s1_req_addr_reg[39]_0 [0]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_req_addr[39]_i_22 
       (.I0(_T_2770[9]),
        .I1(\s1_req_addr_reg[39] [7]),
        .I2(\s1_req_addr_reg[39] [8]),
        .O(\s1_req_addr_reg[39]_1 [3]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_req_addr[39]_i_23 
       (.I0(_T_2770[6]),
        .I1(\s1_req_addr_reg[39] [5]),
        .I2(\s1_req_addr_reg[39] [6]),
        .O(\s1_req_addr_reg[39]_1 [2]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_req_addr[39]_i_24 
       (.I0(\s1_req_addr_reg[39] [2]),
        .I1(\s1_req_addr_reg[39] [3]),
        .I2(\s1_req_addr_reg[39] [4]),
        .O(\s1_req_addr_reg[39]_1 [1]));
  LUT3 #(
    .INIT(8'h01)) 
    \s1_req_addr[39]_i_25 
       (.I0(\s1_req_addr_reg[39] [0]),
        .I1(_T_2770[1]),
        .I2(\s1_req_addr_reg[39] [1]),
        .O(\s1_req_addr_reg[39]_1 [0]));
  LUT1 #(
    .INIT(2'h1)) 
    \s1_req_addr[39]_i_5 
       (.I0(neg_out_reg),
        .O(\s1_req_addr_reg[39] [18]));
  LUT6 #(
    .INIT(64'h00000000C7F7FFFF)) 
    \s1_req_addr[39]_i_7 
       (.I0(_T_2518),
        .I1(ex_reg_rs_lsb_0[1]),
        .I2(ex_reg_rs_lsb_0[0]),
        .I3(_T_2177[24]),
        .I4(ex_reg_rs_bypass_0_reg_0),
        .I5(div_n_526),
        .O(\s1_req_addr_reg[39]_4 ));
  LUT3 #(
    .INIT(8'h80)) 
    \s1_req_addr[39]_i_9 
       (.I0(\s1_req_addr_reg[39] [15]),
        .I1(\s1_req_addr_reg[39] [16]),
        .I2(\s1_req_addr_reg[39] [17]),
        .O(\s1_req_addr_reg[39]_2 [3]));
  (* SOFT_HLUTNM = "soft_lutpair1884" *) 
  LUT2 #(
    .INIT(4'hB)) 
    s1_valid_i_1__1
       (.I0(mem_reg_replay_reg_0),
        .I1(io_mask),
        .O(s1_valid_reg));
  LUT6 #(
    .INIT(64'h0A0A0B0B0B0A0B0A)) 
    s1_valid_i_5
       (.I0(\s1_req_cmd_reg[4] [4]),
        .I1(\s1_req_cmd_reg[4] [3]),
        .I2(\state_reg[0]_1 ),
        .I3(\s1_req_cmd_reg[4] [0]),
        .I4(\s1_req_cmd_reg[4] [2]),
        .I5(\s1_req_cmd_reg[4] [1]),
        .O(\state_reg[1] ));
  (* SOFT_HLUTNM = "soft_lutpair1863" *) 
  LUT2 #(
    .INIT(4'h8)) 
    tag_array_0_reg_i_53
       (.I0(ex_ctrl_mem),
        .I1(ex_reg_valid),
        .O(dcacheArb_io_requestor_1_req_valid));
  (* SOFT_HLUTNM = "soft_lutpair1826" *) 
  LUT5 #(
    .INIT(32'h0020FFEF)) 
    \trig_jalr_count[0]_i_1 
       (.I0(\a_data_reg[63] [0]),
        .I1(\trig_state_reg[0]_0 ),
        .I2(\trig_state_reg[1]_0 ),
        .I3(\trig_state_reg[1]_1 ),
        .I4(trig_jalr_count_reg__0[0]),
        .O(p_0_in__0[0]));
  LUT6 #(
    .INIT(64'hFFEF00200020FFEF)) 
    \trig_jalr_count[1]_i_1 
       (.I0(\a_data_reg[63] [1]),
        .I1(\trig_state_reg[0]_0 ),
        .I2(\trig_state_reg[1]_0 ),
        .I3(\trig_state_reg[1]_1 ),
        .I4(trig_jalr_count_reg__0[0]),
        .I5(trig_jalr_count_reg__0[1]),
        .O(p_0_in__0[1]));
  LUT5 #(
    .INIT(32'hB8B8B88B)) 
    \trig_jalr_count[2]_i_1 
       (.I0(\a_data_reg[63] [2]),
        .I1(\trig_state_reg[0]_1 ),
        .I2(trig_jalr_count_reg__0[2]),
        .I3(trig_jalr_count_reg__0[1]),
        .I4(trig_jalr_count_reg__0[0]),
        .O(p_0_in__0[2]));
  LUT6 #(
    .INIT(64'hB8B8B8B8B8B8B88B)) 
    \trig_jalr_count[3]_i_1 
       (.I0(\a_data_reg[63] [3]),
        .I1(\trig_state_reg[0]_1 ),
        .I2(trig_jalr_count_reg__0[3]),
        .I3(trig_jalr_count_reg__0[2]),
        .I4(trig_jalr_count_reg__0[0]),
        .I5(trig_jalr_count_reg__0[1]),
        .O(p_0_in__0[3]));
  LUT6 #(
    .INIT(64'h00F4004400440044)) 
    \trig_jalr_count[4]_i_1 
       (.I0(\trig_mem_data_reg[127]_0 ),
        .I1(\trig_state_reg[0]_1 ),
        .I2(\trig_jalr_count_reg[0]_0 ),
        .I3(\trig_state_reg[1]_2 ),
        .I4(mem_ctrl_jalr),
        .I5(\trig_jalr_count[4]_i_3_n_0 ),
        .O(trig_jalr_count));
  LUT6 #(
    .INIT(64'h0020FFEFFFEF0020)) 
    \trig_jalr_count[4]_i_2 
       (.I0(\a_data_reg[63] [4]),
        .I1(\trig_state_reg[0]_0 ),
        .I2(\trig_state_reg[1]_0 ),
        .I3(\trig_state_reg[1]_1 ),
        .I4(trig_jalr_count_reg__0[4]),
        .I5(\trig_jalr_count[4]_i_4_n_0 ),
        .O(p_0_in__0[4]));
  (* SOFT_HLUTNM = "soft_lutpair1841" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \trig_jalr_count[4]_i_3 
       (.I0(trig_jalr_count_reg__0[4]),
        .I1(trig_jalr_count_reg__0[3]),
        .I2(trig_jalr_count_reg__0[1]),
        .I3(trig_jalr_count_reg__0[0]),
        .I4(trig_jalr_count_reg__0[2]),
        .O(\trig_jalr_count[4]_i_3_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1841" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \trig_jalr_count[4]_i_4 
       (.I0(trig_jalr_count_reg__0[2]),
        .I1(trig_jalr_count_reg__0[0]),
        .I2(trig_jalr_count_reg__0[1]),
        .I3(trig_jalr_count_reg__0[3]),
        .O(\trig_jalr_count[4]_i_4_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_jalr_count_reg[0] 
       (.C(host_clk),
        .CE(trig_jalr_count),
        .D(p_0_in__0[0]),
        .Q(trig_jalr_count_reg__0[0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_jalr_count_reg[1] 
       (.C(host_clk),
        .CE(trig_jalr_count),
        .D(p_0_in__0[1]),
        .Q(trig_jalr_count_reg__0[1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_jalr_count_reg[2] 
       (.C(host_clk),
        .CE(trig_jalr_count),
        .D(p_0_in__0[2]),
        .Q(trig_jalr_count_reg__0[2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_jalr_count_reg[3] 
       (.C(host_clk),
        .CE(trig_jalr_count),
        .D(p_0_in__0[3]),
        .Q(trig_jalr_count_reg__0[3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_jalr_count_reg[4] 
       (.C(host_clk),
        .CE(trig_jalr_count),
        .D(p_0_in__0[4]),
        .Q(trig_jalr_count_reg__0[4]),
        .R(\<const0> ));
  (* SOFT_HLUTNM = "soft_lutpair1886" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \trig_mem_data[120]_i_1 
       (.I0(\trig_mem_data_reg_n_0_[0] ),
        .I1(_GEN_277[120]),
        .O(\trig_mem_data[120]_i_1_n_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1886" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \trig_mem_data[125]_i_1 
       (.I0(\trig_mem_data_reg_n_0_[0] ),
        .I1(_GEN_277[125]),
        .O(\trig_mem_data[125]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \trig_mem_data[126]_i_1 
       (.I0(\trig_mem_data_reg_n_0_[0] ),
        .I1(\trig_mem_data_reg[126]_0 [1]),
        .O(\trig_mem_data[126]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \trig_mem_data[127]_i_1 
       (.I0(\trig_mem_data[127]_i_2_n_0 ),
        .I1(\trig_mem_data[127]_i_3_n_0 ),
        .I2(\trig_mem_data[127]_i_4_n_0 ),
        .I3(\trig_mem_data[127]_i_5_n_0 ),
        .O(_T_1927));
  LUT5 #(
    .INIT(32'hFFFFFBFF)) 
    \trig_mem_data[127]_i_10 
       (.I0(_GEN_277[24]),
        .I1(_GEN_277[32]),
        .I2(_GEN_277[22]),
        .I3(_GEN_277[52]),
        .I4(\trig_mem_data[127]_i_14_n_0 ),
        .O(\trig_mem_data[127]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hFFDF)) 
    \trig_mem_data[127]_i_11 
       (.I0(_GEN_277[5]),
        .I1(_GEN_277[18]),
        .I2(_GEN_277[51]),
        .I3(_GEN_277[15]),
        .O(\trig_mem_data[127]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF7FF)) 
    \trig_mem_data[127]_i_12 
       (.I0(_GEN_277[0]),
        .I1(_GEN_277[16]),
        .I2(_GEN_277[12]),
        .I3(_GEN_277[9]),
        .I4(\trig_mem_data[127]_i_15_n_0 ),
        .O(\trig_mem_data[127]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \trig_mem_data[127]_i_13 
       (.I0(_GEN_277[45]),
        .I1(_GEN_277[43]),
        .I2(_GEN_277[28]),
        .I3(_GEN_277[3]),
        .O(\trig_mem_data[127]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \trig_mem_data[127]_i_14 
       (.I0(_GEN_277[26]),
        .I1(_GEN_277[11]),
        .I2(_GEN_277[37]),
        .I3(_GEN_277[21]),
        .O(\trig_mem_data[127]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \trig_mem_data[127]_i_15 
       (.I0(_GEN_277[27]),
        .I1(_GEN_277[20]),
        .I2(_GEN_277[31]),
        .I3(_GEN_277[7]),
        .O(\trig_mem_data[127]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBF)) 
    \trig_mem_data[127]_i_2 
       (.I0(\trig_mem_data[127]_i_6_n_0 ),
        .I1(_GEN_277[47]),
        .I2(_GEN_277[40]),
        .I3(_GEN_277[35]),
        .I4(_GEN_277[34]),
        .I5(\trig_mem_data[127]_i_7_n_0 ),
        .O(\trig_mem_data[127]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF7)) 
    \trig_mem_data[127]_i_3 
       (.I0(_GEN_277[13]),
        .I1(_GEN_277[53]),
        .I2(_GEN_277[33]),
        .I3(_GEN_277[36]),
        .I4(\trig_mem_data[127]_i_8_n_0 ),
        .O(\trig_mem_data[127]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \trig_mem_data[127]_i_4 
       (.I0(\trig_mem_data[127]_i_9_n_0 ),
        .I1(_GEN_277[44]),
        .I2(_GEN_277[19]),
        .I3(_GEN_277[6]),
        .I4(_GEN_277[4]),
        .I5(\trig_mem_data[127]_i_10_n_0 ),
        .O(\trig_mem_data[127]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFBFFF)) 
    \trig_mem_data[127]_i_5 
       (.I0(\trig_mem_data[127]_i_11_n_0 ),
        .I1(_GEN_277[25]),
        .I2(\trig_mem_data_reg_n_0_[0] ),
        .I3(_GEN_277[23]),
        .I4(_GEN_277[30]),
        .I5(\trig_mem_data[127]_i_12_n_0 ),
        .O(\trig_mem_data[127]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFFEF)) 
    \trig_mem_data[127]_i_6 
       (.I0(_GEN_277[54]),
        .I1(_GEN_277[8]),
        .I2(_GEN_277[17]),
        .I3(_GEN_277[2]),
        .O(\trig_mem_data[127]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFBFF)) 
    \trig_mem_data[127]_i_7 
       (.I0(_GEN_277[38]),
        .I1(_GEN_277[48]),
        .I2(_GEN_277[1]),
        .I3(_GEN_277[50]),
        .I4(\trig_mem_data[127]_i_13_n_0 ),
        .O(\trig_mem_data[127]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \trig_mem_data[127]_i_8 
       (.I0(_GEN_277[46]),
        .I1(_GEN_277[10]),
        .I2(_GEN_277[49]),
        .I3(_GEN_277[42]),
        .O(\trig_mem_data[127]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \trig_mem_data[127]_i_9 
       (.I0(_GEN_277[39]),
        .I1(_GEN_277[14]),
        .I2(_GEN_277[41]),
        .I3(_GEN_277[29]),
        .O(\trig_mem_data[127]_i_9_n_0 ));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[0] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[0]),
        .Q(\trig_mem_data_reg_n_0_[0] ),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[100] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[100]),
        .Q(_GEN_277[99]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[101] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[101]),
        .Q(_GEN_277[100]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[102] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[102]),
        .Q(_GEN_277[101]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[103] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[103]),
        .Q(_GEN_277[102]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[104] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[104]),
        .Q(_GEN_277[103]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[105] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[105]),
        .Q(_GEN_277[104]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[106] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[106]),
        .Q(_GEN_277[105]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[107] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[107]),
        .Q(_GEN_277[106]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[108] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[108]),
        .Q(_GEN_277[107]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[109] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[109]),
        .Q(_GEN_277[108]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[10] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[10]),
        .Q(_GEN_277[9]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[110] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[110]),
        .Q(_GEN_277[109]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[111] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[111]),
        .Q(_GEN_277[110]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[112] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[112]),
        .Q(_GEN_277[111]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[113] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[113]),
        .Q(_GEN_277[112]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[114] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[114]),
        .Q(_GEN_277[113]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[115] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[115]),
        .Q(_GEN_277[114]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[116] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[116]),
        .Q(_GEN_277[115]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[117] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[117]),
        .Q(_GEN_277[116]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[118] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[118]),
        .Q(_GEN_277[117]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[119] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[119]),
        .Q(_GEN_277[118]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[11] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[11]),
        .Q(_GEN_277[10]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[120] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(\trig_mem_data[120]_i_1_n_0 ),
        .Q(_GEN_277[119]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[121] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[121]),
        .Q(_GEN_277[120]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[122] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[122]),
        .Q(_GEN_277[121]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[123] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[123]),
        .Q(_GEN_277[122]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[124] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[124]),
        .Q(_GEN_277[123]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[125] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(\trig_mem_data[125]_i_1_n_0 ),
        .Q(_GEN_277[124]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[126] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(\trig_mem_data[126]_i_1_n_0 ),
        .Q(_GEN_277[125]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[127] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(\trig_mem_data_reg_n_0_[0] ),
        .Q(\trig_mem_data_reg[126]_0 [1]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[12] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[12]),
        .Q(_GEN_277[11]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[13] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[13]),
        .Q(_GEN_277[12]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[14] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[14]),
        .Q(_GEN_277[13]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[15] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[15]),
        .Q(_GEN_277[14]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[16] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[16]),
        .Q(_GEN_277[15]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[17] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[17]),
        .Q(_GEN_277[16]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[18] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[18]),
        .Q(_GEN_277[17]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[19] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[19]),
        .Q(_GEN_277[18]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[1] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[1]),
        .Q(_GEN_277[0]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[20] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[20]),
        .Q(_GEN_277[19]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[21] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[21]),
        .Q(_GEN_277[20]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[22] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[22]),
        .Q(_GEN_277[21]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[23] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[23]),
        .Q(_GEN_277[22]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[24] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[24]),
        .Q(_GEN_277[23]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[25] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[25]),
        .Q(_GEN_277[24]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[26] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[26]),
        .Q(_GEN_277[25]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[27] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[27]),
        .Q(_GEN_277[26]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[28] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[28]),
        .Q(_GEN_277[27]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[29] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[29]),
        .Q(_GEN_277[28]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[2] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[2]),
        .Q(_GEN_277[1]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[30] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[30]),
        .Q(_GEN_277[29]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[31] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[31]),
        .Q(_GEN_277[30]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[32] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[32]),
        .Q(_GEN_277[31]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[33] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[33]),
        .Q(_GEN_277[32]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[34] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[34]),
        .Q(_GEN_277[33]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[35] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[35]),
        .Q(_GEN_277[34]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[36] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[36]),
        .Q(_GEN_277[35]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[37] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[37]),
        .Q(_GEN_277[36]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[38] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[38]),
        .Q(_GEN_277[37]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[39] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[39]),
        .Q(_GEN_277[38]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[3] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[3]),
        .Q(_GEN_277[2]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[40] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[40]),
        .Q(_GEN_277[39]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[41] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[41]),
        .Q(_GEN_277[40]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[42] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[42]),
        .Q(_GEN_277[41]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[43] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[43]),
        .Q(_GEN_277[42]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[44] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[44]),
        .Q(_GEN_277[43]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[45] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[45]),
        .Q(_GEN_277[44]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[46] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[46]),
        .Q(_GEN_277[45]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[47] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[47]),
        .Q(_GEN_277[46]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[48] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[48]),
        .Q(_GEN_277[47]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[49] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[49]),
        .Q(_GEN_277[48]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[4] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[4]),
        .Q(_GEN_277[3]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[50] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[50]),
        .Q(_GEN_277[49]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[51] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[51]),
        .Q(_GEN_277[50]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[52] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[52]),
        .Q(_GEN_277[51]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[53] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[53]),
        .Q(_GEN_277[52]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[54] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[54]),
        .Q(_GEN_277[53]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[55] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[55]),
        .Q(_GEN_277[54]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[56] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[56]),
        .Q(_GEN_277[55]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[57] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[57]),
        .Q(_GEN_277[56]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[58] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[58]),
        .Q(_GEN_277[57]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[59] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[59]),
        .Q(_GEN_277[58]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[5] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[5]),
        .Q(_GEN_277[4]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[60] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[60]),
        .Q(_GEN_277[59]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[61] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[61]),
        .Q(_GEN_277[60]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[62] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(\trig_mem_data_reg[126]_0 [0]),
        .Q(_GEN_277[61]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[63] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[63]),
        .Q(\trig_mem_data_reg[126]_0 [0]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[64] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[64]),
        .Q(_GEN_277[63]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[65] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[65]),
        .Q(_GEN_277[64]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[66] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[66]),
        .Q(_GEN_277[65]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[67] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[67]),
        .Q(_GEN_277[66]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[68] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[68]),
        .Q(_GEN_277[67]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[69] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[69]),
        .Q(_GEN_277[68]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[6] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[6]),
        .Q(_GEN_277[5]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[70] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[70]),
        .Q(_GEN_277[69]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[71] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[71]),
        .Q(_GEN_277[70]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[72] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[72]),
        .Q(_GEN_277[71]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[73] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[73]),
        .Q(_GEN_277[72]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[74] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[74]),
        .Q(_GEN_277[73]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[75] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[75]),
        .Q(_GEN_277[74]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[76] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[76]),
        .Q(_GEN_277[75]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[77] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[77]),
        .Q(_GEN_277[76]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[78] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[78]),
        .Q(_GEN_277[77]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[79] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[79]),
        .Q(_GEN_277[78]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[7] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[7]),
        .Q(_GEN_277[6]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[80] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[80]),
        .Q(_GEN_277[79]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[81] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[81]),
        .Q(_GEN_277[80]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[82] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[82]),
        .Q(_GEN_277[81]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[83] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[83]),
        .Q(_GEN_277[82]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[84] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[84]),
        .Q(_GEN_277[83]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[85] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[85]),
        .Q(_GEN_277[84]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[86] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[86]),
        .Q(_GEN_277[85]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[87] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[87]),
        .Q(_GEN_277[86]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[88] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[88]),
        .Q(_GEN_277[87]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[89] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[89]),
        .Q(_GEN_277[88]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[8] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[8]),
        .Q(_GEN_277[7]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[90] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[90]),
        .Q(_GEN_277[89]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[91] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[91]),
        .Q(_GEN_277[90]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[92] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[92]),
        .Q(_GEN_277[91]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[93] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[93]),
        .Q(_GEN_277[92]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[94] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[94]),
        .Q(_GEN_277[93]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[95] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[95]),
        .Q(_GEN_277[94]),
        .R(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[96] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[96]),
        .Q(_GEN_277[95]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[97] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[97]),
        .Q(_GEN_277[96]),
        .S(target_reset));
  FDSE #(
    .INIT(1'b1)) 
    \trig_mem_data_reg[98] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[98]),
        .Q(_GEN_277[97]),
        .S(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[99] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[99]),
        .Q(_GEN_277[98]),
        .R(target_reset));
  FDRE #(
    .INIT(1'b0)) 
    \trig_mem_data_reg[9] 
       (.C(host_clk),
        .CE(_T_1927),
        .D(_GEN_277[9]),
        .Q(_GEN_277[8]),
        .R(target_reset));
  LUT6 #(
    .INIT(64'h0000000000040404)) 
    \trig_pc[0]_i_1 
       (.I0(\trig_state_reg[1]_1 ),
        .I1(\trig_state_reg[1]_0 ),
        .I2(\trig_state_reg[0]_0 ),
        .I3(\trig_pc_reg[0]_0 ),
        .I4(\trig_pc_reg[63]_1 ),
        .I5(\trig_mem_data_reg[127]_0 ),
        .O(\trig_pc[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0300010000000100)) 
    \trig_pc[63]_i_1 
       (.I0(\trig_mem_data_reg[127]_0 ),
        .I1(\trig_state_reg[1]_2 ),
        .I2(\trig_state_reg[1]_1 ),
        .I3(\trig_state_reg[1]_0 ),
        .I4(\trig_state_reg[0]_0 ),
        .I5(\trig_pc_reg[0]_1 ),
        .O(trig_pc));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_11 
       (.I0(\a_data_reg[63] [59]),
        .I1(_GEN_277[122]),
        .I2(\a_data_reg[63] [58]),
        .I3(_GEN_277[121]),
        .I4(_GEN_277[120]),
        .I5(\a_data_reg[63] [57]),
        .O(\trig_jalr_count_reg[0]_5 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_12 
       (.I0(_GEN_277[119]),
        .I1(\a_data_reg[63] [56]),
        .I2(\a_data_reg[63] [54]),
        .I3(_GEN_277[117]),
        .I4(\a_data_reg[63] [55]),
        .I5(_GEN_277[118]),
        .O(\trig_jalr_count_reg[0]_5 [2]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_13 
       (.I0(_GEN_277[116]),
        .I1(\a_data_reg[63] [53]),
        .I2(\a_data_reg[63] [51]),
        .I3(_GEN_277[114]),
        .I4(\a_data_reg[63] [52]),
        .I5(_GEN_277[115]),
        .O(\trig_jalr_count_reg[0]_5 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_14 
       (.I0(_GEN_277[113]),
        .I1(\a_data_reg[63] [50]),
        .I2(\a_data_reg[63] [48]),
        .I3(_GEN_277[111]),
        .I4(\a_data_reg[63] [49]),
        .I5(_GEN_277[112]),
        .O(\trig_jalr_count_reg[0]_5 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_16 
       (.I0(_GEN_277[110]),
        .I1(\a_data_reg[63] [47]),
        .I2(\a_data_reg[63] [45]),
        .I3(_GEN_277[108]),
        .I4(\a_data_reg[63] [46]),
        .I5(_GEN_277[109]),
        .O(\trig_jalr_count_reg[0]_4 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_17 
       (.I0(_GEN_277[107]),
        .I1(\a_data_reg[63] [44]),
        .I2(\a_data_reg[63] [42]),
        .I3(_GEN_277[105]),
        .I4(\a_data_reg[63] [43]),
        .I5(_GEN_277[106]),
        .O(\trig_jalr_count_reg[0]_4 [2]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_18 
       (.I0(\a_data_reg[63] [41]),
        .I1(_GEN_277[104]),
        .I2(\a_data_reg[63] [39]),
        .I3(_GEN_277[102]),
        .I4(_GEN_277[103]),
        .I5(\a_data_reg[63] [40]),
        .O(\trig_jalr_count_reg[0]_4 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_19 
       (.I0(_GEN_277[101]),
        .I1(\a_data_reg[63] [38]),
        .I2(\a_data_reg[63] [36]),
        .I3(_GEN_277[99]),
        .I4(\a_data_reg[63] [37]),
        .I5(_GEN_277[100]),
        .O(\trig_jalr_count_reg[0]_4 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_21 
       (.I0(\a_data_reg[63] [35]),
        .I1(_GEN_277[98]),
        .I2(\a_data_reg[63] [33]),
        .I3(_GEN_277[96]),
        .I4(_GEN_277[97]),
        .I5(\a_data_reg[63] [34]),
        .O(\trig_jalr_count_reg[0]_3 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_22 
       (.I0(\a_data_reg[63] [32]),
        .I1(_GEN_277[95]),
        .I2(\a_data_reg[63] [30]),
        .I3(_GEN_277[93]),
        .I4(_GEN_277[94]),
        .I5(\a_data_reg[63] [31]),
        .O(\trig_jalr_count_reg[0]_3 [2]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_23 
       (.I0(\a_data_reg[63] [29]),
        .I1(_GEN_277[92]),
        .I2(\a_data_reg[63] [27]),
        .I3(_GEN_277[90]),
        .I4(_GEN_277[91]),
        .I5(\a_data_reg[63] [28]),
        .O(\trig_jalr_count_reg[0]_3 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_24 
       (.I0(\a_data_reg[63] [24]),
        .I1(_GEN_277[87]),
        .I2(\a_data_reg[63] [25]),
        .I3(_GEN_277[88]),
        .I4(_GEN_277[89]),
        .I5(\a_data_reg[63] [26]),
        .O(\trig_jalr_count_reg[0]_3 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_26 
       (.I0(_GEN_277[86]),
        .I1(\a_data_reg[63] [23]),
        .I2(\a_data_reg[63] [21]),
        .I3(_GEN_277[84]),
        .I4(\a_data_reg[63] [22]),
        .I5(_GEN_277[85]),
        .O(\trig_jalr_count_reg[0]_2 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_27 
       (.I0(_GEN_277[83]),
        .I1(\a_data_reg[63] [20]),
        .I2(\a_data_reg[63] [19]),
        .I3(_GEN_277[82]),
        .I4(\a_data_reg[63] [18]),
        .I5(_GEN_277[81]),
        .O(\trig_jalr_count_reg[0]_2 [2]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_28 
       (.I0(\a_data_reg[63] [17]),
        .I1(_GEN_277[80]),
        .I2(\a_data_reg[63] [15]),
        .I3(_GEN_277[78]),
        .I4(_GEN_277[79]),
        .I5(\a_data_reg[63] [16]),
        .O(\trig_jalr_count_reg[0]_2 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_29 
       (.I0(\a_data_reg[63] [14]),
        .I1(_GEN_277[77]),
        .I2(\a_data_reg[63] [12]),
        .I3(_GEN_277[75]),
        .I4(_GEN_277[76]),
        .I5(\a_data_reg[63] [13]),
        .O(\trig_jalr_count_reg[0]_2 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_30 
       (.I0(_GEN_277[73]),
        .I1(\a_data_reg[63] [10]),
        .I2(\a_data_reg[63] [11]),
        .I3(_GEN_277[74]),
        .I4(\a_data_reg[63] [9]),
        .I5(_GEN_277[72]),
        .O(\trig_jalr_count_reg[0]_1 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_31 
       (.I0(_GEN_277[71]),
        .I1(\a_data_reg[63] [8]),
        .I2(\a_data_reg[63] [7]),
        .I3(_GEN_277[70]),
        .I4(\a_data_reg[63] [6]),
        .I5(_GEN_277[69]),
        .O(\trig_jalr_count_reg[0]_1 [2]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_32 
       (.I0(_GEN_277[68]),
        .I1(\a_data_reg[63] [5]),
        .I2(\a_data_reg[63] [4]),
        .I3(_GEN_277[67]),
        .I4(\a_data_reg[63] [3]),
        .I5(_GEN_277[66]),
        .O(\trig_jalr_count_reg[0]_1 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_33 
       (.I0(_GEN_277[65]),
        .I1(\a_data_reg[63] [2]),
        .I2(\a_data_reg[63] [0]),
        .I3(_GEN_277[63]),
        .I4(\a_data_reg[63] [1]),
        .I5(_GEN_277[64]),
        .O(\trig_jalr_count_reg[0]_1 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_pc[63]_i_9 
       (.I0(\a_data_reg[63] [62]),
        .I1(_GEN_277[125]),
        .I2(\a_data_reg[63] [60]),
        .I3(_GEN_277[123]),
        .I4(_GEN_277[124]),
        .I5(\a_data_reg[63] [61]),
        .O(\trig_jalr_count_reg[0]_6 ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[0] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[0]),
        .Q(\trig_pc_reg[63]_0 [0]),
        .R(\trig_pc[0]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[10] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[10]),
        .Q(\trig_pc_reg[63]_0 [10]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[11] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[11]),
        .Q(\trig_pc_reg[63]_0 [11]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[12] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[12]),
        .Q(\trig_pc_reg[63]_0 [12]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[13] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[13]),
        .Q(\trig_pc_reg[63]_0 [13]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[14] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[14]),
        .Q(\trig_pc_reg[63]_0 [14]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[15] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[15]),
        .Q(\trig_pc_reg[63]_0 [15]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[16] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[16]),
        .Q(\trig_pc_reg[63]_0 [16]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[17] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[17]),
        .Q(\trig_pc_reg[63]_0 [17]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[18] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[18]),
        .Q(\trig_pc_reg[63]_0 [18]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[19] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[19]),
        .Q(\trig_pc_reg[63]_0 [19]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[1] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[1]),
        .Q(\trig_pc_reg[63]_0 [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[20] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[20]),
        .Q(\trig_pc_reg[63]_0 [20]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[21] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[21]),
        .Q(\trig_pc_reg[63]_0 [21]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[22] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[22]),
        .Q(\trig_pc_reg[63]_0 [22]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[23] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[23]),
        .Q(\trig_pc_reg[63]_0 [23]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[24] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[24]),
        .Q(\trig_pc_reg[63]_0 [24]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[25] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[25]),
        .Q(\trig_pc_reg[63]_0 [25]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[26] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[26]),
        .Q(\trig_pc_reg[63]_0 [26]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[27] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[27]),
        .Q(\trig_pc_reg[63]_0 [27]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[28] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[28]),
        .Q(\trig_pc_reg[63]_0 [28]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[29] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[29]),
        .Q(\trig_pc_reg[63]_0 [29]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[2] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[2]),
        .Q(\trig_pc_reg[63]_0 [2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[30] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[30]),
        .Q(\trig_pc_reg[63]_0 [30]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[31] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[31]),
        .Q(\trig_pc_reg[63]_0 [31]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[32] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[32]),
        .Q(\trig_pc_reg[63]_0 [32]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[33] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[33]),
        .Q(\trig_pc_reg[63]_0 [33]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[34] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[34]),
        .Q(\trig_pc_reg[63]_0 [34]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[35] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[35]),
        .Q(\trig_pc_reg[63]_0 [35]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[36] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[36]),
        .Q(\trig_pc_reg[63]_0 [36]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[37] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[37]),
        .Q(\trig_pc_reg[63]_0 [37]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[38] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[38]),
        .Q(\trig_pc_reg[63]_0 [38]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[39] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[39]),
        .Q(\trig_pc_reg[63]_0 [39]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[3] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[3]),
        .Q(\trig_pc_reg[63]_0 [3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[40] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[40]),
        .Q(\trig_pc_reg[63]_0 [40]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[41] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[41]),
        .Q(\trig_pc_reg[63]_0 [41]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[42] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[42]),
        .Q(\trig_pc_reg[63]_0 [42]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[43] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[43]),
        .Q(\trig_pc_reg[63]_0 [43]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[44] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[44]),
        .Q(\trig_pc_reg[63]_0 [44]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[45] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[45]),
        .Q(\trig_pc_reg[63]_0 [45]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[46] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[46]),
        .Q(\trig_pc_reg[63]_0 [46]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[47] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[47]),
        .Q(\trig_pc_reg[63]_0 [47]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[48] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[48]),
        .Q(\trig_pc_reg[63]_0 [48]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[49] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[49]),
        .Q(\trig_pc_reg[63]_0 [49]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[4] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[4]),
        .Q(\trig_pc_reg[63]_0 [4]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[50] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[50]),
        .Q(\trig_pc_reg[63]_0 [50]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[51] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[51]),
        .Q(\trig_pc_reg[63]_0 [51]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[52] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[52]),
        .Q(\trig_pc_reg[63]_0 [52]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[53] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[53]),
        .Q(\trig_pc_reg[63]_0 [53]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[54] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[54]),
        .Q(\trig_pc_reg[63]_0 [54]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[55] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[55]),
        .Q(\trig_pc_reg[63]_0 [55]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[56] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[56]),
        .Q(\trig_pc_reg[63]_0 [56]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[57] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[57]),
        .Q(\trig_pc_reg[63]_0 [57]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[58] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[58]),
        .Q(\trig_pc_reg[63]_0 [58]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[59] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[59]),
        .Q(\trig_pc_reg[63]_0 [59]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[5] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[5]),
        .Q(\trig_pc_reg[63]_0 [5]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[60] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[60]),
        .Q(\trig_pc_reg[63]_0 [60]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[61] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[61]),
        .Q(\trig_pc_reg[63]_0 [61]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[62] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[62]),
        .Q(\trig_pc_reg[63]_0 [62]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[63] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[63]),
        .Q(\trig_pc_reg[63]_0 [63]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[6] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[6]),
        .Q(\trig_pc_reg[63]_0 [6]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[7] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[7]),
        .Q(\trig_pc_reg[63]_0 [7]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[8] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[8]),
        .Q(\trig_pc_reg[63]_0 [8]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_pc_reg[9] 
       (.C(host_clk),
        .CE(trig_pc),
        .D(out[9]),
        .Q(\trig_pc_reg[63]_0 [9]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    trig_pc_valid_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(trig_pc_valid_reg_1),
        .Q(\trig_pc_reg[0]_0 ),
        .R(target_reset));
  LUT6 #(
    .INIT(64'h0000000000E2E2E2)) 
    \trig_state[0]_i_1 
       (.I0(\trig_state_reg[0]_0 ),
        .I1(\trig_state[0]_i_2_n_0 ),
        .I2(trig_state),
        .I3(\trig_state[0]_i_4_n_0 ),
        .I4(\trig_state_reg[1]_2 ),
        .I5(target_reset),
        .O(\trig_state[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00AA00FF00FF88F0)) 
    \trig_state[0]_i_2 
       (.I0(trig_pc_valid_reg_2),
        .I1(mem_ctrl_branch),
        .I2(\trig_mem_data_reg[63]_0 ),
        .I3(\trig_state_reg[1]_1 ),
        .I4(\trig_state_reg[0]_0 ),
        .I5(\trig_state_reg[1]_0 ),
        .O(\trig_state[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000C5F)) 
    \trig_state[0]_i_3 
       (.I0(\trig_mem_data_reg[127]_0 ),
        .I1(\trig_mem_data_reg[63]_0 ),
        .I2(\trig_state_reg[1]_0 ),
        .I3(\trig_state_reg[0]_0 ),
        .I4(\trig_state_reg[1]_1 ),
        .I5(\trig_state_reg[1]_2 ),
        .O(trig_state));
  LUT3 #(
    .INIT(8'h01)) 
    \trig_state[0]_i_4 
       (.I0(\trig_state_reg[1]_1 ),
        .I1(\trig_state_reg[0]_0 ),
        .I2(\trig_state_reg[1]_0 ),
        .O(\trig_state[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000A8A8A8AA)) 
    \trig_state[1]_i_1 
       (.I0(\trig_state[1]_i_2_n_0 ),
        .I1(\trig_state_reg[1]_1 ),
        .I2(\trig_state_reg[1]_0 ),
        .I3(\trig_state_reg[1]_2 ),
        .I4(\trig_mem_data_reg[63]_0 ),
        .I5(target_reset),
        .O(\trig_state[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_10 
       (.I0(_GEN_277[52]),
        .I1(\a_data_reg[63] [53]),
        .I2(\a_data_reg[63] [51]),
        .I3(_GEN_277[50]),
        .I4(\a_data_reg[63] [52]),
        .I5(_GEN_277[51]),
        .O(\trig_state_reg[1]_7 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_11 
       (.I0(_GEN_277[49]),
        .I1(\a_data_reg[63] [50]),
        .I2(\a_data_reg[63] [48]),
        .I3(_GEN_277[47]),
        .I4(\a_data_reg[63] [49]),
        .I5(_GEN_277[48]),
        .O(\trig_state_reg[1]_7 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_13 
       (.I0(_GEN_277[46]),
        .I1(\a_data_reg[63] [47]),
        .I2(\a_data_reg[63] [45]),
        .I3(_GEN_277[44]),
        .I4(\a_data_reg[63] [46]),
        .I5(_GEN_277[45]),
        .O(\trig_state_reg[1]_6 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_14 
       (.I0(_GEN_277[43]),
        .I1(\a_data_reg[63] [44]),
        .I2(\a_data_reg[63] [43]),
        .I3(_GEN_277[42]),
        .I4(\a_data_reg[63] [42]),
        .I5(_GEN_277[41]),
        .O(\trig_state_reg[1]_6 [2]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_15 
       (.I0(\a_data_reg[63] [39]),
        .I1(_GEN_277[38]),
        .I2(\a_data_reg[63] [40]),
        .I3(_GEN_277[39]),
        .I4(_GEN_277[40]),
        .I5(\a_data_reg[63] [41]),
        .O(\trig_state_reg[1]_6 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_16 
       (.I0(_GEN_277[37]),
        .I1(\a_data_reg[63] [38]),
        .I2(\a_data_reg[63] [36]),
        .I3(_GEN_277[35]),
        .I4(\a_data_reg[63] [37]),
        .I5(_GEN_277[36]),
        .O(\trig_state_reg[1]_6 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_18 
       (.I0(\a_data_reg[63] [33]),
        .I1(_GEN_277[32]),
        .I2(\a_data_reg[63] [34]),
        .I3(_GEN_277[33]),
        .I4(_GEN_277[34]),
        .I5(\a_data_reg[63] [35]),
        .O(\trig_state_reg[1]_5 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_19 
       (.I0(\a_data_reg[63] [30]),
        .I1(_GEN_277[29]),
        .I2(\a_data_reg[63] [31]),
        .I3(_GEN_277[30]),
        .I4(_GEN_277[31]),
        .I5(\a_data_reg[63] [32]),
        .O(\trig_state_reg[1]_5 [2]));
  LUT6 #(
    .INIT(64'h0101FFFF04000000)) 
    \trig_state[1]_i_2 
       (.I0(\trig_state_reg[1]_2 ),
        .I1(\trig_state_reg[0]_0 ),
        .I2(\trig_state_reg[1]_1 ),
        .I3(\trig_mem_data_reg[127]_0 ),
        .I4(\trig_state[1]_i_4_n_0 ),
        .I5(\trig_state_reg[1]_0 ),
        .O(\trig_state[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_20 
       (.I0(\a_data_reg[63] [28]),
        .I1(_GEN_277[27]),
        .I2(\a_data_reg[63] [27]),
        .I3(_GEN_277[26]),
        .I4(_GEN_277[28]),
        .I5(\a_data_reg[63] [29]),
        .O(\trig_state_reg[1]_5 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_21 
       (.I0(\a_data_reg[63] [26]),
        .I1(_GEN_277[25]),
        .I2(\a_data_reg[63] [24]),
        .I3(_GEN_277[23]),
        .I4(_GEN_277[24]),
        .I5(\a_data_reg[63] [25]),
        .O(\trig_state_reg[1]_5 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_23 
       (.I0(_GEN_277[22]),
        .I1(\a_data_reg[63] [23]),
        .I2(\a_data_reg[63] [21]),
        .I3(_GEN_277[20]),
        .I4(\a_data_reg[63] [22]),
        .I5(_GEN_277[21]),
        .O(\trig_state_reg[1]_4 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_24 
       (.I0(_GEN_277[19]),
        .I1(\a_data_reg[63] [20]),
        .I2(\a_data_reg[63] [18]),
        .I3(_GEN_277[17]),
        .I4(\a_data_reg[63] [19]),
        .I5(_GEN_277[18]),
        .O(\trig_state_reg[1]_4 [2]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_25 
       (.I0(\a_data_reg[63] [15]),
        .I1(_GEN_277[14]),
        .I2(\a_data_reg[63] [16]),
        .I3(_GEN_277[15]),
        .I4(_GEN_277[16]),
        .I5(\a_data_reg[63] [17]),
        .O(\trig_state_reg[1]_4 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_26 
       (.I0(\a_data_reg[63] [12]),
        .I1(_GEN_277[11]),
        .I2(\a_data_reg[63] [13]),
        .I3(_GEN_277[12]),
        .I4(_GEN_277[13]),
        .I5(\a_data_reg[63] [14]),
        .O(\trig_state_reg[1]_4 [0]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_27 
       (.I0(_GEN_277[9]),
        .I1(\a_data_reg[63] [10]),
        .I2(\a_data_reg[63] [11]),
        .I3(_GEN_277[10]),
        .I4(\a_data_reg[63] [9]),
        .I5(_GEN_277[8]),
        .O(\trig_state_reg[1]_3 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_28 
       (.I0(_GEN_277[7]),
        .I1(\a_data_reg[63] [8]),
        .I2(\a_data_reg[63] [6]),
        .I3(_GEN_277[5]),
        .I4(\a_data_reg[63] [7]),
        .I5(_GEN_277[6]),
        .O(\trig_state_reg[1]_3 [2]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_29 
       (.I0(_GEN_277[4]),
        .I1(\a_data_reg[63] [5]),
        .I2(\a_data_reg[63] [3]),
        .I3(_GEN_277[2]),
        .I4(\a_data_reg[63] [4]),
        .I5(_GEN_277[3]),
        .O(\trig_state_reg[1]_3 [1]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_30 
       (.I0(_GEN_277[1]),
        .I1(\a_data_reg[63] [2]),
        .I2(\a_data_reg[63] [1]),
        .I3(_GEN_277[0]),
        .I4(\a_data_reg[63] [0]),
        .I5(\trig_mem_data_reg_n_0_[0] ),
        .O(\trig_state_reg[1]_3 [0]));
  LUT6 #(
    .INIT(64'h000FEFF00000EFF0)) 
    \trig_state[1]_i_4 
       (.I0(\trig_pc_reg[0]_1 ),
        .I1(\trig_state_reg[1]_2 ),
        .I2(\trig_state_reg[0]_0 ),
        .I3(\trig_state_reg[1]_0 ),
        .I4(\trig_state_reg[1]_1 ),
        .I5(mem_ctrl_branch),
        .O(\trig_state[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_6 
       (.I0(\a_data_reg[63] [60]),
        .I1(_GEN_277[59]),
        .I2(\a_data_reg[63] [61]),
        .I3(_GEN_277[60]),
        .I4(_GEN_277[61]),
        .I5(\a_data_reg[63] [62]),
        .O(\trig_state_reg[1]_8 ));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_8 
       (.I0(\a_data_reg[63] [59]),
        .I1(_GEN_277[58]),
        .I2(\a_data_reg[63] [57]),
        .I3(_GEN_277[56]),
        .I4(_GEN_277[57]),
        .I5(\a_data_reg[63] [58]),
        .O(\trig_state_reg[1]_7 [3]));
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \trig_state[1]_i_9 
       (.I0(_GEN_277[55]),
        .I1(\a_data_reg[63] [56]),
        .I2(\a_data_reg[63] [54]),
        .I3(_GEN_277[53]),
        .I4(\a_data_reg[63] [55]),
        .I5(_GEN_277[54]),
        .O(\trig_state_reg[1]_7 [2]));
  FDRE #(
    .INIT(1'b0)) 
    \trig_state_reg[0] 
       (.C(host_clk),
        .CE(\<const1> ),
        .D(\trig_state[0]_i_1_n_0 ),
        .Q(\trig_state_reg[0]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_state_reg[1] 
       (.C(host_clk),
        .CE(\<const1> ),
        .D(\trig_state[1]_i_1_n_0 ),
        .Q(\trig_state_reg[1]_0 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \trig_state_reg[2] 
       (.C(host_clk),
        .CE(\<const1> ),
        .D(mem_ctrl_branch_reg_0),
        .Q(\trig_state_reg[1]_1 ),
        .R(target_reset));
  (* SOFT_HLUTNM = "soft_lutpair1879" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \valid[3]_i_3__0 
       (.I0(frontend_io_cpu_sfence_valid),
        .I1(s2_replay),
        .O(\valid_reg[3] ));
  LUT6 #(
    .INIT(64'hEEEEEEEEEEEEEEFE)) 
    \valid[4]_i_1__0 
       (.I0(p_2_in),
        .I1(target_reset),
        .I2(frontend_io_cpu_sfence_valid),
        .I3(s2_replay),
        .I4(frontend_io_cpu_sfence_bits_rs2),
        .I5(\valid_reg[3]_1 ),
        .O(\valid_reg[3]_0 ));
  (* SOFT_HLUTNM = "soft_lutpair1849" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \valid[4]_i_4 
       (.I0(wb_reg_valid),
        .I1(wb_reg_sfence),
        .O(frontend_io_cpu_sfence_valid));
  (* SOFT_HLUTNM = "soft_lutpair1849" *) 
  LUT4 #(
    .INIT(16'hFF08)) 
    \vb_array[63]_i_1 
       (.I0(wb_ctrl_fence_i),
        .I1(wb_reg_valid),
        .I2(dcacheArb_io_requestor_1_s2_nack),
        .I3(target_reset),
        .O(SR));
  FDRE #(
    .INIT(1'b0)) 
    \wb_ctrl_csr_reg[0] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_ctrl_csr[0]),
        .Q(\reg_sscratch_reg[59] [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_ctrl_csr_reg[1] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_ctrl_csr[1]),
        .Q(\reg_sscratch_reg[59] [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_ctrl_csr_reg[2] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_ctrl_csr[2]),
        .Q(\reg_sscratch_reg[59] [2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    wb_ctrl_div_reg
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_ctrl_div),
        .Q(wb_ctrl_div),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    wb_ctrl_fence_i_reg
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(wb_ctrl_fence_i_reg_0),
        .Q(wb_ctrl_fence_i),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'hFE)) 
    wb_ctrl_mem_i_1
       (.I0(mem_reg_replay),
        .I1(mem_reg_xcpt_interrupt),
        .I2(mem_reg_valid),
        .O(mem_pc_valid));
  FDRE #(
    .INIT(1'b0)) 
    wb_ctrl_mem_reg
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_ctrl_mem),
        .Q(wb_ctrl_mem),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_ctrl_mem_type_reg[0] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\mem_ctrl_mem_type_reg_n_0_[0] ),
        .Q(\valid_reg[3]_1 ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_ctrl_mem_type_reg[1] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\mem_ctrl_mem_type_reg_n_0_[1] ),
        .Q(frontend_io_cpu_sfence_bits_rs2),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    wb_ctrl_wxd_reg
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_ctrl_wxd),
        .Q(wb_ctrl_wxd),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'hA8)) 
    \wb_reg_cause[63]_i_1 
       (.I0(mem_reg_cause[63]),
        .I1(mem_reg_xcpt),
        .I2(mem_reg_xcpt_interrupt),
        .O(\wb_reg_cause[63]_i_1_n_0 ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_cause_reg[0] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(csr_n_748),
        .Q(wb_reg_cause[0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_cause_reg[1] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(csr_n_747),
        .Q(wb_reg_cause[1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_cause_reg[2] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_reg_xcpt_interrupt_reg_0[0]),
        .Q(\reg_scause_reg[2] ),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_cause_reg[3] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_reg_xcpt_interrupt_reg_0[1]),
        .Q(wb_reg_cause[3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_cause_reg[63] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_cause[63]_i_1_n_0 ),
        .Q(wb_reg_cause[63]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    wb_reg_flush_pipe_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(wb_reg_flush_pipe0),
        .Q(wb_reg_flush_pipe),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[10] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [3]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[11] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [4]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [4]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[20] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [13]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [5]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[21] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [14]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [6]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[22] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [15]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [7]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[23] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [16]),
        .Q(csr_io_rw_addr[3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[24] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [17]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [8]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[25] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [18]),
        .Q(csr_io_rw_addr[5]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[26] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [19]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [9]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[27] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [20]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [10]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[28] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [21]),
        .Q(csr_io_rw_addr[8]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[29] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [22]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [11]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[30] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [23]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [12]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[31] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [24]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [13]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[7] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [0]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[8] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [1]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_inst_reg[9] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_inst_reg[31]_0 [2]),
        .Q(\reg_bp_0_control_tmatch_reg[1] [2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[10] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [9]),
        .Q(\reg_dpc_reg[39] [9]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[11] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [10]),
        .Q(\reg_dpc_reg[39] [10]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[12] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [11]),
        .Q(\reg_dpc_reg[39] [11]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[13] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [12]),
        .Q(\reg_dpc_reg[39] [12]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[14] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [13]),
        .Q(\reg_dpc_reg[39] [13]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[15] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [14]),
        .Q(\reg_dpc_reg[39] [14]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[16] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [15]),
        .Q(\reg_dpc_reg[39] [15]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[17] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [16]),
        .Q(\reg_dpc_reg[39] [16]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[18] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [17]),
        .Q(\reg_dpc_reg[39] [17]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[19] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [18]),
        .Q(\reg_dpc_reg[39] [18]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[1] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [0]),
        .Q(\reg_dpc_reg[39] [0]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[20] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [19]),
        .Q(\reg_dpc_reg[39] [19]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[21] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [20]),
        .Q(\reg_dpc_reg[39] [20]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[22] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [21]),
        .Q(\reg_dpc_reg[39] [21]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[23] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [22]),
        .Q(\reg_dpc_reg[39] [22]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[24] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [23]),
        .Q(\reg_dpc_reg[39] [23]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[25] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [24]),
        .Q(\reg_dpc_reg[39] [24]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[26] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [25]),
        .Q(\reg_dpc_reg[39] [25]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[27] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [26]),
        .Q(\reg_dpc_reg[39] [26]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[28] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\bypass_mux_2_reg[31]_0 [0]),
        .Q(\reg_dpc_reg[39] [27]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[29] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\bypass_mux_2_reg[31]_0 [1]),
        .Q(\reg_dpc_reg[39] [28]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[2] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [1]),
        .Q(\reg_dpc_reg[39] [1]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[30] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\bypass_mux_2_reg[31]_0 [2]),
        .Q(\reg_dpc_reg[39] [29]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[31] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [27]),
        .Q(\reg_dpc_reg[39] [30]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[32] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[34]_0 [1]),
        .Q(\reg_dpc_reg[39] [31]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[33] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[34]_0 [2]),
        .Q(\reg_dpc_reg[39] [32]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[34] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[34]_0 [3]),
        .Q(\reg_dpc_reg[39] [33]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[35] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [28]),
        .Q(\reg_dpc_reg[39] [34]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[36] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [29]),
        .Q(\reg_dpc_reg[39] [35]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[37] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [30]),
        .Q(\reg_dpc_reg[39] [36]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[38] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [31]),
        .Q(\reg_dpc_reg[39] [37]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[39] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [32]),
        .Q(\reg_dpc_reg[39] [38]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[3] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [2]),
        .Q(\reg_dpc_reg[39] [2]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[4] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [3]),
        .Q(\reg_dpc_reg[39] [3]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[5] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [4]),
        .Q(\reg_dpc_reg[39] [4]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[6] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [5]),
        .Q(\reg_dpc_reg[39] [5]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[7] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [6]),
        .Q(\reg_dpc_reg[39] [6]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[8] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [7]),
        .Q(\reg_dpc_reg[39] [7]),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    \wb_reg_pc_reg[9] 
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(\wb_reg_pc_reg[39]_0 [8]),
        .Q(\reg_dpc_reg[39] [8]),
        .R(\<const0> ));
  LUT5 #(
    .INIT(32'hAAAA8000)) 
    wb_reg_replay_i_1
       (.I0(frontend_io_cpu_req_bits_speculative),
        .I1(dcacheArb_io_requestor_1_replay_next),
        .I2(mem_ctrl_wxd),
        .I3(mem_reg_valid),
        .I4(mem_reg_replay),
        .O(wb_reg_replay0));
  FDRE #(
    .INIT(1'b0)) 
    wb_reg_replay_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(wb_reg_replay0),
        .Q(wb_reg_replay),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    wb_reg_sfence_reg
       (.C(host_clk),
        .CE(mem_pc_valid),
        .D(mem_reg_sfence),
        .Q(wb_reg_sfence),
        .R(\<const0> ));
  FDRE #(
    .INIT(1'b0)) 
    wb_reg_valid_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(_T_2377),
        .Q(wb_reg_valid),
        .R(\<const0> ));
  LUT5 #(
    .INIT(32'h0000FFEA)) 
    wb_reg_xcpt_i_2
       (.I0(\reg_bp_0_control_tmatch_reg[1] [7]),
        .I1(\reg_bp_0_control_tmatch_reg[1] [5]),
        .I2(\reg_bp_0_control_tmatch_reg[1] [6]),
        .I3(\wb_ctrl_csr_reg[0]_0 ),
        .I4(dcache_io_cpu_invalidate_lr),
        .O(wb_reg_xcpt_i_2_n_0));
  FDRE #(
    .INIT(1'b0)) 
    wb_reg_xcpt_reg
       (.C(host_clk),
        .CE(\<const1> ),
        .D(wb_reg_xcpt0),
        .Q(wb_reg_xcpt),
        .R(\<const0> ));
endmodule 